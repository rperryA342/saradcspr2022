magic
tech sky130A
timestamp 1649877290
<< metal3 >>
rect 710 805 810 905
rect -220 -225 810 805
<< mimcap >>
rect -205 689 795 790
rect -205 589 -106 689
rect -6 589 69 689
rect 169 589 244 689
rect 344 589 419 689
rect 519 589 594 689
rect 694 589 795 689
rect -205 514 795 589
rect -205 414 -106 514
rect -6 414 69 514
rect 169 414 244 514
rect 344 414 419 514
rect 519 414 594 514
rect 694 414 795 514
rect -205 339 795 414
rect -205 239 -106 339
rect -6 239 69 339
rect 169 239 244 339
rect 344 239 419 339
rect 519 239 594 339
rect 694 239 795 339
rect -205 164 795 239
rect -205 64 -106 164
rect -6 64 69 164
rect 169 64 244 164
rect 344 64 419 164
rect 519 64 594 164
rect 694 64 795 164
rect -205 -11 795 64
rect -205 -111 -106 -11
rect -6 -111 69 -11
rect 169 -111 244 -11
rect 344 -111 419 -11
rect 519 -111 594 -11
rect 694 -111 795 -11
rect -205 -210 795 -111
<< mimcapcontact >>
rect -106 589 -6 689
rect 69 589 169 689
rect 244 589 344 689
rect 419 589 519 689
rect 594 589 694 689
rect -106 414 -6 514
rect 69 414 169 514
rect 244 414 344 514
rect 419 414 519 514
rect 594 414 694 514
rect -106 239 -6 339
rect 69 239 169 339
rect 244 239 344 339
rect 419 239 519 339
rect 594 239 694 339
rect -106 64 -6 164
rect 69 64 169 164
rect 244 64 344 164
rect 419 64 519 164
rect 594 64 694 164
rect -106 -111 -6 -11
rect 69 -111 169 -11
rect 244 -111 344 -11
rect 419 -111 519 -11
rect 594 -111 694 -11
<< metal4 >>
rect 207 739 383 740
rect -156 689 744 739
rect -156 589 -106 689
rect -6 589 69 689
rect 169 589 244 689
rect 344 589 419 689
rect 519 589 594 689
rect 694 589 744 689
rect -156 514 744 589
rect -156 414 -106 514
rect -6 414 69 514
rect 169 414 244 514
rect 344 414 419 514
rect 519 414 594 514
rect 694 414 744 514
rect -156 339 744 414
rect -156 239 -106 339
rect -6 239 69 339
rect 169 239 244 339
rect 344 239 419 339
rect 519 239 594 339
rect 694 239 744 339
rect -156 164 744 239
rect -156 64 -106 164
rect -6 64 69 164
rect 169 64 244 164
rect 344 64 419 164
rect 519 64 594 164
rect 694 64 744 164
rect -156 -11 744 64
rect -156 -111 -106 -11
rect -6 -111 69 -11
rect 169 -111 244 -11
rect 344 -111 419 -11
rect 519 -111 594 -11
rect 694 -111 744 -11
rect -156 -160 744 -111
rect -156 -161 205 -160
rect 245 -375 345 -160
rect 385 -161 744 -160
<< labels >>
rlabel metal4 295 -375 295 -375 5 top1C
rlabel metal3 765 905 765 905 1 common
<< end >>
