magic
tech sky130A
magscale 1 2
timestamp 1651353626
<< checkpaint >>
rect -3932 -3932 18676 20820
<< viali >>
rect 1501 14569 1535 14603
rect 6653 14569 6687 14603
rect 10517 14569 10551 14603
rect 12817 14569 12851 14603
rect 1685 14365 1719 14399
rect 2697 14365 2731 14399
rect 6837 14365 6871 14399
rect 10701 14365 10735 14399
rect 12633 14365 12667 14399
rect 2881 14229 2915 14263
rect 6377 13889 6411 13923
rect 9413 13889 9447 13923
rect 10241 13889 10275 13923
rect 10057 13821 10091 13855
rect 4261 13685 4295 13719
rect 6561 13685 6595 13719
rect 9229 13685 9263 13719
rect 10701 13481 10735 13515
rect 4261 13345 4295 13379
rect 6837 13345 6871 13379
rect 9229 13345 9263 13379
rect 3893 13277 3927 13311
rect 6561 13277 6595 13311
rect 8953 13277 8987 13311
rect 12633 13277 12667 13311
rect 5687 13141 5721 13175
rect 8309 13141 8343 13175
rect 12817 13141 12851 13175
rect 6837 12937 6871 12971
rect 9689 12937 9723 12971
rect 10057 12937 10091 12971
rect 4997 12801 5031 12835
rect 5089 12801 5123 12835
rect 5273 12801 5307 12835
rect 5365 12801 5399 12835
rect 6377 12801 6411 12835
rect 12357 12801 12391 12835
rect 10149 12733 10183 12767
rect 10241 12733 10275 12767
rect 6653 12665 6687 12699
rect 12173 12665 12207 12699
rect 4813 12597 4847 12631
rect 6377 12393 6411 12427
rect 4629 12257 4663 12291
rect 4905 12257 4939 12291
rect 9597 12189 9631 12223
rect 9873 12121 9907 12155
rect 11345 12053 11379 12087
rect 9781 11849 9815 11883
rect 2697 11781 2731 11815
rect 1685 11713 1719 11747
rect 6929 11713 6963 11747
rect 2421 11645 2455 11679
rect 4169 11645 4203 11679
rect 8033 11645 8067 11679
rect 8309 11645 8343 11679
rect 1501 11577 1535 11611
rect 7113 11577 7147 11611
rect 8401 11305 8435 11339
rect 12817 11305 12851 11339
rect 6653 11169 6687 11203
rect 11069 11169 11103 11203
rect 11345 11169 11379 11203
rect 3985 11101 4019 11135
rect 4261 11101 4295 11135
rect 4445 11101 4479 11135
rect 9505 11101 9539 11135
rect 6929 11033 6963 11067
rect 9321 11033 9355 11067
rect 3801 10965 3835 10999
rect 2053 10761 2087 10795
rect 3525 10693 3559 10727
rect 8125 10693 8159 10727
rect 8677 10625 8711 10659
rect 8861 10625 8895 10659
rect 9137 10625 9171 10659
rect 9965 10625 9999 10659
rect 10241 10625 10275 10659
rect 10425 10625 10459 10659
rect 3801 10557 3835 10591
rect 9321 10557 9355 10591
rect 8033 10421 8067 10455
rect 9781 10421 9815 10455
rect 7665 10217 7699 10251
rect 9781 10081 9815 10115
rect 11253 10081 11287 10115
rect 12725 10081 12759 10115
rect 4077 10013 4111 10047
rect 4353 10013 4387 10047
rect 4537 10013 4571 10047
rect 4997 10013 5031 10047
rect 5917 10013 5951 10047
rect 9505 10013 9539 10047
rect 12449 10013 12483 10047
rect 6193 9945 6227 9979
rect 3893 9877 3927 9911
rect 5181 9877 5215 9911
rect 12081 9877 12115 9911
rect 12541 9877 12575 9911
rect 4261 9605 4295 9639
rect 6745 9605 6779 9639
rect 6929 9537 6963 9571
rect 9229 9537 9263 9571
rect 12173 9537 12207 9571
rect 1501 9469 1535 9503
rect 1777 9469 1811 9503
rect 3249 9469 3283 9503
rect 3985 9469 4019 9503
rect 9045 9469 9079 9503
rect 9137 9469 9171 9503
rect 9597 9401 9631 9435
rect 5733 9333 5767 9367
rect 11989 9333 12023 9367
rect 2605 9129 2639 9163
rect 6745 9129 6779 9163
rect 12909 9129 12943 9163
rect 3801 9061 3835 9095
rect 4445 8993 4479 9027
rect 5273 8993 5307 9027
rect 11437 8993 11471 9027
rect 2789 8925 2823 8959
rect 3065 8925 3099 8959
rect 3249 8925 3283 8959
rect 4997 8925 5031 8959
rect 11161 8925 11195 8959
rect 4169 8857 4203 8891
rect 4261 8789 4295 8823
rect 4169 8585 4203 8619
rect 9597 8585 9631 8619
rect 12817 8585 12851 8619
rect 3985 8449 4019 8483
rect 9413 8449 9447 8483
rect 12633 8449 12667 8483
rect 11161 8041 11195 8075
rect 9229 7905 9263 7939
rect 12909 7905 12943 7939
rect 1685 7837 1719 7871
rect 2329 7837 2363 7871
rect 3801 7837 3835 7871
rect 6837 7837 6871 7871
rect 7113 7837 7147 7871
rect 7297 7837 7331 7871
rect 7941 7837 7975 7871
rect 8217 7837 8251 7871
rect 8401 7837 8435 7871
rect 8953 7837 8987 7871
rect 7757 7769 7791 7803
rect 12633 7769 12667 7803
rect 1501 7701 1535 7735
rect 2145 7701 2179 7735
rect 3985 7701 4019 7735
rect 6653 7701 6687 7735
rect 10701 7701 10735 7735
rect 3157 7497 3191 7531
rect 8585 7497 8619 7531
rect 10977 7497 11011 7531
rect 12725 7497 12759 7531
rect 1685 7429 1719 7463
rect 6653 7429 6687 7463
rect 3617 7361 3651 7395
rect 4445 7361 4479 7395
rect 8769 7361 8803 7395
rect 12081 7361 12115 7395
rect 12817 7361 12851 7395
rect 1409 7293 1443 7327
rect 6377 7293 6411 7327
rect 9229 7293 9263 7327
rect 9505 7293 9539 7327
rect 3801 7225 3835 7259
rect 4261 7157 4295 7191
rect 8125 7157 8159 7191
rect 11989 7157 12023 7191
rect 2329 6953 2363 6987
rect 4242 6953 4276 6987
rect 6929 6953 6963 6987
rect 2881 6817 2915 6851
rect 3985 6817 4019 6851
rect 7573 6817 7607 6851
rect 9229 6817 9263 6851
rect 10517 6817 10551 6851
rect 10793 6817 10827 6851
rect 12265 6817 12299 6851
rect 2697 6749 2731 6783
rect 7297 6749 7331 6783
rect 9505 6749 9539 6783
rect 2789 6613 2823 6647
rect 5733 6613 5767 6647
rect 7389 6613 7423 6647
rect 3157 6409 3191 6443
rect 7205 6409 7239 6443
rect 7297 6341 7331 6375
rect 4905 6273 4939 6307
rect 4629 6205 4663 6239
rect 12817 5797 12851 5831
rect 4537 5729 4571 5763
rect 9689 5729 9723 5763
rect 9965 5661 9999 5695
rect 11069 5661 11103 5695
rect 11345 5661 11379 5695
rect 11529 5661 11563 5695
rect 4261 5593 4295 5627
rect 12633 5593 12667 5627
rect 3893 5525 3927 5559
rect 4353 5525 4387 5559
rect 9873 5525 9907 5559
rect 10333 5525 10367 5559
rect 10885 5525 10919 5559
rect 3893 5321 3927 5355
rect 10057 5321 10091 5355
rect 7481 5253 7515 5287
rect 4077 5185 4111 5219
rect 4353 5185 4387 5219
rect 4537 5185 4571 5219
rect 5181 5185 5215 5219
rect 5457 5185 5491 5219
rect 5641 5185 5675 5219
rect 9413 5185 9447 5219
rect 9597 5185 9631 5219
rect 9873 5185 9907 5219
rect 10701 5185 10735 5219
rect 12633 5185 12667 5219
rect 4997 5117 5031 5151
rect 7205 5117 7239 5151
rect 8953 5117 8987 5151
rect 12909 5117 12943 5151
rect 10609 4981 10643 5015
rect 6469 4641 6503 4675
rect 8953 4641 8987 4675
rect 9229 4641 9263 4675
rect 11437 4641 11471 4675
rect 2145 4573 2179 4607
rect 3801 4573 3835 4607
rect 11161 4573 11195 4607
rect 6193 4505 6227 4539
rect 2329 4437 2363 4471
rect 3985 4437 4019 4471
rect 4721 4437 4755 4471
rect 10701 4437 10735 4471
rect 12909 4437 12943 4471
rect 2697 4233 2731 4267
rect 4997 4233 5031 4267
rect 9229 4233 9263 4267
rect 12725 4233 12759 4267
rect 6929 4165 6963 4199
rect 10701 4165 10735 4199
rect 2329 4097 2363 4131
rect 3249 4097 3283 4131
rect 7021 4097 7055 4131
rect 8125 4097 8159 4131
rect 8309 4097 8343 4131
rect 8585 4097 8619 4131
rect 10977 4097 11011 4131
rect 12909 4097 12943 4131
rect 2145 4029 2179 4063
rect 2237 4029 2271 4063
rect 3525 4029 3559 4063
rect 7113 4029 7147 4063
rect 6561 3893 6595 3927
rect 8769 3893 8803 3927
rect 1409 3689 1443 3723
rect 3985 3689 4019 3723
rect 7573 3689 7607 3723
rect 8401 3689 8435 3723
rect 10701 3689 10735 3723
rect 2881 3553 2915 3587
rect 9229 3553 9263 3587
rect 3157 3485 3191 3519
rect 3801 3485 3835 3519
rect 5825 3485 5859 3519
rect 8217 3485 8251 3519
rect 8953 3485 8987 3519
rect 6101 3417 6135 3451
rect 1501 3145 1535 3179
rect 2421 3145 2455 3179
rect 6377 3145 6411 3179
rect 7021 3077 7055 3111
rect 7205 3077 7239 3111
rect 1685 3009 1719 3043
rect 4169 3009 4203 3043
rect 6561 3009 6595 3043
rect 3893 2941 3927 2975
rect 3249 2601 3283 2635
rect 2053 2533 2087 2567
rect 4353 2465 4387 2499
rect 3065 2397 3099 2431
rect 4077 2397 4111 2431
rect 7849 2397 7883 2431
rect 11713 2397 11747 2431
rect 12633 2397 12667 2431
rect 1869 2329 1903 2363
rect 8033 2261 8067 2295
rect 11897 2261 11931 2295
rect 12817 2261 12851 2295
<< metal1 >>
rect 1104 14714 13616 14736
rect 1104 14662 2514 14714
rect 2566 14662 2578 14714
rect 2630 14662 2642 14714
rect 2694 14662 2706 14714
rect 2758 14662 2770 14714
rect 2822 14662 5642 14714
rect 5694 14662 5706 14714
rect 5758 14662 5770 14714
rect 5822 14662 5834 14714
rect 5886 14662 5898 14714
rect 5950 14662 8770 14714
rect 8822 14662 8834 14714
rect 8886 14662 8898 14714
rect 8950 14662 8962 14714
rect 9014 14662 9026 14714
rect 9078 14662 11898 14714
rect 11950 14662 11962 14714
rect 12014 14662 12026 14714
rect 12078 14662 12090 14714
rect 12142 14662 12154 14714
rect 12206 14662 13616 14714
rect 1104 14640 13616 14662
rect 1486 14600 1492 14612
rect 1447 14572 1492 14600
rect 1486 14560 1492 14572
rect 1544 14560 1550 14612
rect 6454 14560 6460 14612
rect 6512 14600 6518 14612
rect 6641 14603 6699 14609
rect 6641 14600 6653 14603
rect 6512 14572 6653 14600
rect 6512 14560 6518 14572
rect 6641 14569 6653 14572
rect 6687 14569 6699 14603
rect 6641 14563 6699 14569
rect 10318 14560 10324 14612
rect 10376 14600 10382 14612
rect 10505 14603 10563 14609
rect 10505 14600 10517 14603
rect 10376 14572 10517 14600
rect 10376 14560 10382 14572
rect 10505 14569 10517 14572
rect 10551 14569 10563 14603
rect 10505 14563 10563 14569
rect 12805 14603 12863 14609
rect 12805 14569 12817 14603
rect 12851 14600 12863 14603
rect 14182 14600 14188 14612
rect 12851 14572 14188 14600
rect 12851 14569 12863 14572
rect 12805 14563 12863 14569
rect 14182 14560 14188 14572
rect 14240 14560 14246 14612
rect 1673 14399 1731 14405
rect 1673 14365 1685 14399
rect 1719 14365 1731 14399
rect 1673 14359 1731 14365
rect 1688 14328 1716 14359
rect 2406 14356 2412 14408
rect 2464 14396 2470 14408
rect 2685 14399 2743 14405
rect 2685 14396 2697 14399
rect 2464 14368 2697 14396
rect 2464 14356 2470 14368
rect 2685 14365 2697 14368
rect 2731 14365 2743 14399
rect 2685 14359 2743 14365
rect 6825 14399 6883 14405
rect 6825 14365 6837 14399
rect 6871 14396 6883 14399
rect 7006 14396 7012 14408
rect 6871 14368 7012 14396
rect 6871 14365 6883 14368
rect 6825 14359 6883 14365
rect 7006 14356 7012 14368
rect 7064 14356 7070 14408
rect 10686 14396 10692 14408
rect 10647 14368 10692 14396
rect 10686 14356 10692 14368
rect 10744 14356 10750 14408
rect 12434 14356 12440 14408
rect 12492 14396 12498 14408
rect 12621 14399 12679 14405
rect 12621 14396 12633 14399
rect 12492 14368 12633 14396
rect 12492 14356 12498 14368
rect 12621 14365 12633 14368
rect 12667 14365 12679 14399
rect 12621 14359 12679 14365
rect 3234 14328 3240 14340
rect 1688 14300 3240 14328
rect 3234 14288 3240 14300
rect 3292 14288 3298 14340
rect 2869 14263 2927 14269
rect 2869 14229 2881 14263
rect 2915 14260 2927 14263
rect 4982 14260 4988 14272
rect 2915 14232 4988 14260
rect 2915 14229 2927 14232
rect 2869 14223 2927 14229
rect 4982 14220 4988 14232
rect 5040 14220 5046 14272
rect 1104 14170 13616 14192
rect 1104 14118 4078 14170
rect 4130 14118 4142 14170
rect 4194 14118 4206 14170
rect 4258 14118 4270 14170
rect 4322 14118 4334 14170
rect 4386 14118 7206 14170
rect 7258 14118 7270 14170
rect 7322 14118 7334 14170
rect 7386 14118 7398 14170
rect 7450 14118 7462 14170
rect 7514 14118 10334 14170
rect 10386 14118 10398 14170
rect 10450 14118 10462 14170
rect 10514 14118 10526 14170
rect 10578 14118 10590 14170
rect 10642 14118 13616 14170
rect 1104 14096 13616 14118
rect 6362 13920 6368 13932
rect 6323 13892 6368 13920
rect 6362 13880 6368 13892
rect 6420 13880 6426 13932
rect 9401 13923 9459 13929
rect 9401 13889 9413 13923
rect 9447 13920 9459 13923
rect 9766 13920 9772 13932
rect 9447 13892 9772 13920
rect 9447 13889 9459 13892
rect 9401 13883 9459 13889
rect 9766 13880 9772 13892
rect 9824 13880 9830 13932
rect 10226 13920 10232 13932
rect 10187 13892 10232 13920
rect 10226 13880 10232 13892
rect 10284 13880 10290 13932
rect 10042 13852 10048 13864
rect 10003 13824 10048 13852
rect 10042 13812 10048 13824
rect 10100 13812 10106 13864
rect 4246 13716 4252 13728
rect 4207 13688 4252 13716
rect 4246 13676 4252 13688
rect 4304 13676 4310 13728
rect 6549 13719 6607 13725
rect 6549 13685 6561 13719
rect 6595 13716 6607 13719
rect 6822 13716 6828 13728
rect 6595 13688 6828 13716
rect 6595 13685 6607 13688
rect 6549 13679 6607 13685
rect 6822 13676 6828 13688
rect 6880 13676 6886 13728
rect 9214 13716 9220 13728
rect 9175 13688 9220 13716
rect 9214 13676 9220 13688
rect 9272 13676 9278 13728
rect 1104 13626 13616 13648
rect 1104 13574 2514 13626
rect 2566 13574 2578 13626
rect 2630 13574 2642 13626
rect 2694 13574 2706 13626
rect 2758 13574 2770 13626
rect 2822 13574 5642 13626
rect 5694 13574 5706 13626
rect 5758 13574 5770 13626
rect 5822 13574 5834 13626
rect 5886 13574 5898 13626
rect 5950 13574 8770 13626
rect 8822 13574 8834 13626
rect 8886 13574 8898 13626
rect 8950 13574 8962 13626
rect 9014 13574 9026 13626
rect 9078 13574 11898 13626
rect 11950 13574 11962 13626
rect 12014 13574 12026 13626
rect 12078 13574 12090 13626
rect 12142 13574 12154 13626
rect 12206 13574 13616 13626
rect 1104 13552 13616 13574
rect 10686 13512 10692 13524
rect 10647 13484 10692 13512
rect 10686 13472 10692 13484
rect 10744 13472 10750 13524
rect 4246 13376 4252 13388
rect 4207 13348 4252 13376
rect 4246 13336 4252 13348
rect 4304 13336 4310 13388
rect 6822 13376 6828 13388
rect 6783 13348 6828 13376
rect 6822 13336 6828 13348
rect 6880 13336 6886 13388
rect 9214 13376 9220 13388
rect 9175 13348 9220 13376
rect 9214 13336 9220 13348
rect 9272 13336 9278 13388
rect 3881 13311 3939 13317
rect 3881 13277 3893 13311
rect 3927 13308 3939 13311
rect 4338 13308 4344 13320
rect 3927 13280 4344 13308
rect 3927 13277 3939 13280
rect 3881 13271 3939 13277
rect 4338 13268 4344 13280
rect 4396 13268 4402 13320
rect 6546 13308 6552 13320
rect 6507 13280 6552 13308
rect 6546 13268 6552 13280
rect 6604 13268 6610 13320
rect 8941 13311 8999 13317
rect 8941 13277 8953 13311
rect 8987 13277 8999 13311
rect 8941 13271 8999 13277
rect 12621 13311 12679 13317
rect 12621 13277 12633 13311
rect 12667 13308 12679 13311
rect 12986 13308 12992 13320
rect 12667 13280 12992 13308
rect 12667 13277 12679 13280
rect 12621 13271 12679 13277
rect 8202 13240 8208 13252
rect 5290 13212 6914 13240
rect 8050 13212 8208 13240
rect 5442 13132 5448 13184
rect 5500 13172 5506 13184
rect 5675 13175 5733 13181
rect 5675 13172 5687 13175
rect 5500 13144 5687 13172
rect 5500 13132 5506 13144
rect 5675 13141 5687 13144
rect 5721 13141 5733 13175
rect 6886 13172 6914 13212
rect 8128 13172 8156 13212
rect 8202 13200 8208 13212
rect 8260 13200 8266 13252
rect 8956 13240 8984 13271
rect 12986 13268 12992 13280
rect 13044 13268 13050 13320
rect 10962 13240 10968 13252
rect 8956 13212 9628 13240
rect 10442 13212 10968 13240
rect 9600 13184 9628 13212
rect 10962 13200 10968 13212
rect 11020 13200 11026 13252
rect 8294 13172 8300 13184
rect 6886 13144 8156 13172
rect 8255 13144 8300 13172
rect 5675 13135 5733 13141
rect 8294 13132 8300 13144
rect 8352 13132 8358 13184
rect 9582 13132 9588 13184
rect 9640 13132 9646 13184
rect 12802 13172 12808 13184
rect 12763 13144 12808 13172
rect 12802 13132 12808 13144
rect 12860 13132 12866 13184
rect 1104 13082 13616 13104
rect 1104 13030 4078 13082
rect 4130 13030 4142 13082
rect 4194 13030 4206 13082
rect 4258 13030 4270 13082
rect 4322 13030 4334 13082
rect 4386 13030 7206 13082
rect 7258 13030 7270 13082
rect 7322 13030 7334 13082
rect 7386 13030 7398 13082
rect 7450 13030 7462 13082
rect 7514 13030 10334 13082
rect 10386 13030 10398 13082
rect 10450 13030 10462 13082
rect 10514 13030 10526 13082
rect 10578 13030 10590 13082
rect 10642 13030 13616 13082
rect 1104 13008 13616 13030
rect 6362 12928 6368 12980
rect 6420 12968 6426 12980
rect 6825 12971 6883 12977
rect 6825 12968 6837 12971
rect 6420 12940 6837 12968
rect 6420 12928 6426 12940
rect 6825 12937 6837 12940
rect 6871 12937 6883 12971
rect 6825 12931 6883 12937
rect 9677 12971 9735 12977
rect 9677 12937 9689 12971
rect 9723 12968 9735 12971
rect 9766 12968 9772 12980
rect 9723 12940 9772 12968
rect 9723 12937 9735 12940
rect 9677 12931 9735 12937
rect 9766 12928 9772 12940
rect 9824 12928 9830 12980
rect 10045 12971 10103 12977
rect 10045 12937 10057 12971
rect 10091 12968 10103 12971
rect 10686 12968 10692 12980
rect 10091 12940 10692 12968
rect 10091 12937 10103 12940
rect 10045 12931 10103 12937
rect 10686 12928 10692 12940
rect 10744 12928 10750 12980
rect 5000 12872 6408 12900
rect 5000 12844 5028 12872
rect 4982 12832 4988 12844
rect 4943 12804 4988 12832
rect 4982 12792 4988 12804
rect 5040 12792 5046 12844
rect 5077 12835 5135 12841
rect 5077 12801 5089 12835
rect 5123 12801 5135 12835
rect 5258 12832 5264 12844
rect 5219 12804 5264 12832
rect 5077 12795 5135 12801
rect 5092 12696 5120 12795
rect 5258 12792 5264 12804
rect 5316 12792 5322 12844
rect 5353 12835 5411 12841
rect 5353 12801 5365 12835
rect 5399 12832 5411 12835
rect 5442 12832 5448 12844
rect 5399 12804 5448 12832
rect 5399 12801 5411 12804
rect 5353 12795 5411 12801
rect 5442 12792 5448 12804
rect 5500 12792 5506 12844
rect 6380 12841 6408 12872
rect 6365 12835 6423 12841
rect 6365 12801 6377 12835
rect 6411 12801 6423 12835
rect 6365 12795 6423 12801
rect 12345 12835 12403 12841
rect 12345 12801 12357 12835
rect 12391 12832 12403 12835
rect 12710 12832 12716 12844
rect 12391 12804 12716 12832
rect 12391 12801 12403 12804
rect 12345 12795 12403 12801
rect 12710 12792 12716 12804
rect 12768 12792 12774 12844
rect 10134 12764 10140 12776
rect 10095 12736 10140 12764
rect 10134 12724 10140 12736
rect 10192 12724 10198 12776
rect 10226 12724 10232 12776
rect 10284 12764 10290 12776
rect 12802 12764 12808 12776
rect 10284 12736 12808 12764
rect 10284 12724 10290 12736
rect 12802 12724 12808 12736
rect 12860 12724 12866 12776
rect 6270 12696 6276 12708
rect 5092 12668 6276 12696
rect 6270 12656 6276 12668
rect 6328 12696 6334 12708
rect 6641 12699 6699 12705
rect 6641 12696 6653 12699
rect 6328 12668 6653 12696
rect 6328 12656 6334 12668
rect 6641 12665 6653 12668
rect 6687 12665 6699 12699
rect 6641 12659 6699 12665
rect 10962 12656 10968 12708
rect 11020 12696 11026 12708
rect 12161 12699 12219 12705
rect 12161 12696 12173 12699
rect 11020 12668 12173 12696
rect 11020 12656 11026 12668
rect 12161 12665 12173 12668
rect 12207 12665 12219 12699
rect 12161 12659 12219 12665
rect 4801 12631 4859 12637
rect 4801 12597 4813 12631
rect 4847 12628 4859 12631
rect 4890 12628 4896 12640
rect 4847 12600 4896 12628
rect 4847 12597 4859 12600
rect 4801 12591 4859 12597
rect 4890 12588 4896 12600
rect 4948 12588 4954 12640
rect 1104 12538 13616 12560
rect 1104 12486 2514 12538
rect 2566 12486 2578 12538
rect 2630 12486 2642 12538
rect 2694 12486 2706 12538
rect 2758 12486 2770 12538
rect 2822 12486 5642 12538
rect 5694 12486 5706 12538
rect 5758 12486 5770 12538
rect 5822 12486 5834 12538
rect 5886 12486 5898 12538
rect 5950 12486 8770 12538
rect 8822 12486 8834 12538
rect 8886 12486 8898 12538
rect 8950 12486 8962 12538
rect 9014 12486 9026 12538
rect 9078 12486 11898 12538
rect 11950 12486 11962 12538
rect 12014 12486 12026 12538
rect 12078 12486 12090 12538
rect 12142 12486 12154 12538
rect 12206 12486 13616 12538
rect 1104 12464 13616 12486
rect 6270 12384 6276 12436
rect 6328 12424 6334 12436
rect 6365 12427 6423 12433
rect 6365 12424 6377 12427
rect 6328 12396 6377 12424
rect 6328 12384 6334 12396
rect 6365 12393 6377 12396
rect 6411 12393 6423 12427
rect 6365 12387 6423 12393
rect 4430 12248 4436 12300
rect 4488 12288 4494 12300
rect 4614 12288 4620 12300
rect 4488 12260 4620 12288
rect 4488 12248 4494 12260
rect 4614 12248 4620 12260
rect 4672 12248 4678 12300
rect 4890 12288 4896 12300
rect 4851 12260 4896 12288
rect 4890 12248 4896 12260
rect 4948 12248 4954 12300
rect 9582 12220 9588 12232
rect 9543 12192 9588 12220
rect 9582 12180 9588 12192
rect 9640 12180 9646 12232
rect 10962 12180 10968 12232
rect 11020 12180 11026 12232
rect 8202 12152 8208 12164
rect 6118 12124 8208 12152
rect 8202 12112 8208 12124
rect 8260 12112 8266 12164
rect 9122 12112 9128 12164
rect 9180 12152 9186 12164
rect 9861 12155 9919 12161
rect 9861 12152 9873 12155
rect 9180 12124 9873 12152
rect 9180 12112 9186 12124
rect 9861 12121 9873 12124
rect 9907 12121 9919 12155
rect 9861 12115 9919 12121
rect 7926 12044 7932 12096
rect 7984 12084 7990 12096
rect 10042 12084 10048 12096
rect 7984 12056 10048 12084
rect 7984 12044 7990 12056
rect 10042 12044 10048 12056
rect 10100 12044 10106 12096
rect 11330 12084 11336 12096
rect 11291 12056 11336 12084
rect 11330 12044 11336 12056
rect 11388 12044 11394 12096
rect 1104 11994 13616 12016
rect 1104 11942 4078 11994
rect 4130 11942 4142 11994
rect 4194 11942 4206 11994
rect 4258 11942 4270 11994
rect 4322 11942 4334 11994
rect 4386 11942 7206 11994
rect 7258 11942 7270 11994
rect 7322 11942 7334 11994
rect 7386 11942 7398 11994
rect 7450 11942 7462 11994
rect 7514 11942 10334 11994
rect 10386 11942 10398 11994
rect 10450 11942 10462 11994
rect 10514 11942 10526 11994
rect 10578 11942 10590 11994
rect 10642 11942 13616 11994
rect 1104 11920 13616 11942
rect 9122 11840 9128 11892
rect 9180 11880 9186 11892
rect 9769 11883 9827 11889
rect 9769 11880 9781 11883
rect 9180 11852 9781 11880
rect 9180 11840 9186 11852
rect 9769 11849 9781 11852
rect 9815 11849 9827 11883
rect 9769 11843 9827 11849
rect 2406 11772 2412 11824
rect 2464 11812 2470 11824
rect 2685 11815 2743 11821
rect 2685 11812 2697 11815
rect 2464 11784 2697 11812
rect 2464 11772 2470 11784
rect 2685 11781 2697 11784
rect 2731 11781 2743 11815
rect 2685 11775 2743 11781
rect 2958 11772 2964 11824
rect 3016 11812 3022 11824
rect 9674 11812 9680 11824
rect 3016 11784 3174 11812
rect 9522 11784 9680 11812
rect 3016 11772 3022 11784
rect 9674 11772 9680 11784
rect 9732 11812 9738 11824
rect 10962 11812 10968 11824
rect 9732 11784 10968 11812
rect 9732 11772 9738 11784
rect 10962 11772 10968 11784
rect 11020 11772 11026 11824
rect 1673 11747 1731 11753
rect 1673 11713 1685 11747
rect 1719 11744 1731 11747
rect 2038 11744 2044 11756
rect 1719 11716 2044 11744
rect 1719 11713 1731 11716
rect 1673 11707 1731 11713
rect 2038 11704 2044 11716
rect 2096 11704 2102 11756
rect 6546 11704 6552 11756
rect 6604 11744 6610 11756
rect 6917 11747 6975 11753
rect 6917 11744 6929 11747
rect 6604 11716 6929 11744
rect 6604 11704 6610 11716
rect 6917 11713 6929 11716
rect 6963 11713 6975 11747
rect 6917 11707 6975 11713
rect 2314 11636 2320 11688
rect 2372 11676 2378 11688
rect 2409 11679 2467 11685
rect 2409 11676 2421 11679
rect 2372 11648 2421 11676
rect 2372 11636 2378 11648
rect 2409 11645 2421 11648
rect 2455 11645 2467 11679
rect 4154 11676 4160 11688
rect 4067 11648 4160 11676
rect 2409 11639 2467 11645
rect 4154 11636 4160 11648
rect 4212 11676 4218 11688
rect 5258 11676 5264 11688
rect 4212 11648 5264 11676
rect 4212 11636 4218 11648
rect 5258 11636 5264 11648
rect 5316 11636 5322 11688
rect 8021 11679 8079 11685
rect 8021 11645 8033 11679
rect 8067 11645 8079 11679
rect 8021 11639 8079 11645
rect 8297 11679 8355 11685
rect 8297 11645 8309 11679
rect 8343 11676 8355 11679
rect 8386 11676 8392 11688
rect 8343 11648 8392 11676
rect 8343 11645 8355 11648
rect 8297 11639 8355 11645
rect 1486 11608 1492 11620
rect 1447 11580 1492 11608
rect 1486 11568 1492 11580
rect 1544 11568 1550 11620
rect 7101 11611 7159 11617
rect 7101 11577 7113 11611
rect 7147 11608 7159 11611
rect 8036 11608 8064 11639
rect 8386 11636 8392 11648
rect 8444 11636 8450 11688
rect 7147 11580 8064 11608
rect 7147 11577 7159 11580
rect 7101 11571 7159 11577
rect 2406 11500 2412 11552
rect 2464 11540 2470 11552
rect 7926 11540 7932 11552
rect 2464 11512 7932 11540
rect 2464 11500 2470 11512
rect 7926 11500 7932 11512
rect 7984 11500 7990 11552
rect 8036 11540 8064 11580
rect 9582 11540 9588 11552
rect 8036 11512 9588 11540
rect 9582 11500 9588 11512
rect 9640 11500 9646 11552
rect 1104 11450 13616 11472
rect 1104 11398 2514 11450
rect 2566 11398 2578 11450
rect 2630 11398 2642 11450
rect 2694 11398 2706 11450
rect 2758 11398 2770 11450
rect 2822 11398 5642 11450
rect 5694 11398 5706 11450
rect 5758 11398 5770 11450
rect 5822 11398 5834 11450
rect 5886 11398 5898 11450
rect 5950 11398 8770 11450
rect 8822 11398 8834 11450
rect 8886 11398 8898 11450
rect 8950 11398 8962 11450
rect 9014 11398 9026 11450
rect 9078 11398 11898 11450
rect 11950 11398 11962 11450
rect 12014 11398 12026 11450
rect 12078 11398 12090 11450
rect 12142 11398 12154 11450
rect 12206 11398 13616 11450
rect 1104 11376 13616 11398
rect 8386 11336 8392 11348
rect 8347 11308 8392 11336
rect 8386 11296 8392 11308
rect 8444 11296 8450 11348
rect 12802 11336 12808 11348
rect 12763 11308 12808 11336
rect 12802 11296 12808 11308
rect 12860 11296 12866 11348
rect 6546 11160 6552 11212
rect 6604 11200 6610 11212
rect 6641 11203 6699 11209
rect 6641 11200 6653 11203
rect 6604 11172 6653 11200
rect 6604 11160 6610 11172
rect 6641 11169 6653 11172
rect 6687 11169 6699 11203
rect 6641 11163 6699 11169
rect 9582 11160 9588 11212
rect 9640 11200 9646 11212
rect 11057 11203 11115 11209
rect 11057 11200 11069 11203
rect 9640 11172 11069 11200
rect 9640 11160 9646 11172
rect 11057 11169 11069 11172
rect 11103 11169 11115 11203
rect 11330 11200 11336 11212
rect 11291 11172 11336 11200
rect 11057 11163 11115 11169
rect 11330 11160 11336 11172
rect 11388 11160 11394 11212
rect 3973 11135 4031 11141
rect 3973 11101 3985 11135
rect 4019 11132 4031 11135
rect 4154 11132 4160 11144
rect 4019 11104 4160 11132
rect 4019 11101 4031 11104
rect 3973 11095 4031 11101
rect 4154 11092 4160 11104
rect 4212 11092 4218 11144
rect 4249 11135 4307 11141
rect 4249 11101 4261 11135
rect 4295 11101 4307 11135
rect 4430 11132 4436 11144
rect 4391 11104 4436 11132
rect 4249 11095 4307 11101
rect 2038 11024 2044 11076
rect 2096 11064 2102 11076
rect 4264 11064 4292 11095
rect 4430 11092 4436 11104
rect 4488 11092 4494 11144
rect 9493 11135 9551 11141
rect 9493 11101 9505 11135
rect 9539 11132 9551 11135
rect 9674 11132 9680 11144
rect 9539 11104 9680 11132
rect 9539 11101 9551 11104
rect 9493 11095 9551 11101
rect 9674 11092 9680 11104
rect 9732 11092 9738 11144
rect 2096 11036 4292 11064
rect 2096 11024 2102 11036
rect 6914 11024 6920 11076
rect 6972 11064 6978 11076
rect 8202 11064 8208 11076
rect 6972 11036 7017 11064
rect 8115 11036 8208 11064
rect 6972 11024 6978 11036
rect 8202 11024 8208 11036
rect 8260 11064 8266 11076
rect 9309 11067 9367 11073
rect 9309 11064 9321 11067
rect 8260 11036 9321 11064
rect 8260 11024 8266 11036
rect 9309 11033 9321 11036
rect 9355 11033 9367 11067
rect 12710 11064 12716 11076
rect 12558 11036 12716 11064
rect 9309 11027 9367 11033
rect 12710 11024 12716 11036
rect 12768 11024 12774 11076
rect 3786 10996 3792 11008
rect 3747 10968 3792 10996
rect 3786 10956 3792 10968
rect 3844 10956 3850 11008
rect 1104 10906 13616 10928
rect 1104 10854 4078 10906
rect 4130 10854 4142 10906
rect 4194 10854 4206 10906
rect 4258 10854 4270 10906
rect 4322 10854 4334 10906
rect 4386 10854 7206 10906
rect 7258 10854 7270 10906
rect 7322 10854 7334 10906
rect 7386 10854 7398 10906
rect 7450 10854 7462 10906
rect 7514 10854 10334 10906
rect 10386 10854 10398 10906
rect 10450 10854 10462 10906
rect 10514 10854 10526 10906
rect 10578 10854 10590 10906
rect 10642 10854 13616 10906
rect 1104 10832 13616 10854
rect 2038 10792 2044 10804
rect 1999 10764 2044 10792
rect 2038 10752 2044 10764
rect 2096 10752 2102 10804
rect 2866 10684 2872 10736
rect 2924 10684 2930 10736
rect 3513 10727 3571 10733
rect 3513 10693 3525 10727
rect 3559 10724 3571 10727
rect 3786 10724 3792 10736
rect 3559 10696 3792 10724
rect 3559 10693 3571 10696
rect 3513 10687 3571 10693
rect 3786 10684 3792 10696
rect 3844 10684 3850 10736
rect 8113 10727 8171 10733
rect 8113 10693 8125 10727
rect 8159 10724 8171 10727
rect 8294 10724 8300 10736
rect 8159 10696 8300 10724
rect 8159 10693 8171 10696
rect 8113 10687 8171 10693
rect 8294 10684 8300 10696
rect 8352 10684 8358 10736
rect 10134 10684 10140 10736
rect 10192 10724 10198 10736
rect 10192 10696 10456 10724
rect 10192 10684 10198 10696
rect 8312 10656 8340 10684
rect 10428 10668 10456 10696
rect 8665 10659 8723 10665
rect 8665 10656 8677 10659
rect 8312 10628 8677 10656
rect 8665 10625 8677 10628
rect 8711 10625 8723 10659
rect 8665 10619 8723 10625
rect 8849 10659 8907 10665
rect 8849 10625 8861 10659
rect 8895 10625 8907 10659
rect 9122 10656 9128 10668
rect 9083 10628 9128 10656
rect 8849 10619 8907 10625
rect 1394 10548 1400 10600
rect 1452 10588 1458 10600
rect 2314 10588 2320 10600
rect 1452 10560 2320 10588
rect 1452 10548 1458 10560
rect 2314 10548 2320 10560
rect 2372 10588 2378 10600
rect 3789 10591 3847 10597
rect 3789 10588 3801 10591
rect 2372 10560 3801 10588
rect 2372 10548 2378 10560
rect 3789 10557 3801 10560
rect 3835 10557 3847 10591
rect 3789 10551 3847 10557
rect 7650 10548 7656 10600
rect 7708 10588 7714 10600
rect 8864 10588 8892 10619
rect 9122 10616 9128 10628
rect 9180 10616 9186 10668
rect 9950 10656 9956 10668
rect 9911 10628 9956 10656
rect 9950 10616 9956 10628
rect 10008 10616 10014 10668
rect 10229 10659 10287 10665
rect 10229 10625 10241 10659
rect 10275 10625 10287 10659
rect 10410 10656 10416 10668
rect 10371 10628 10416 10656
rect 10229 10619 10287 10625
rect 7708 10560 8892 10588
rect 9309 10591 9367 10597
rect 7708 10548 7714 10560
rect 9309 10557 9321 10591
rect 9355 10588 9367 10591
rect 10244 10588 10272 10619
rect 10410 10616 10416 10628
rect 10468 10616 10474 10668
rect 9355 10560 10272 10588
rect 9355 10557 9367 10560
rect 9309 10551 9367 10557
rect 8021 10455 8079 10461
rect 8021 10421 8033 10455
rect 8067 10452 8079 10455
rect 8110 10452 8116 10464
rect 8067 10424 8116 10452
rect 8067 10421 8079 10424
rect 8021 10415 8079 10421
rect 8110 10412 8116 10424
rect 8168 10412 8174 10464
rect 9766 10452 9772 10464
rect 9727 10424 9772 10452
rect 9766 10412 9772 10424
rect 9824 10412 9830 10464
rect 1104 10362 13616 10384
rect 1104 10310 2514 10362
rect 2566 10310 2578 10362
rect 2630 10310 2642 10362
rect 2694 10310 2706 10362
rect 2758 10310 2770 10362
rect 2822 10310 5642 10362
rect 5694 10310 5706 10362
rect 5758 10310 5770 10362
rect 5822 10310 5834 10362
rect 5886 10310 5898 10362
rect 5950 10310 8770 10362
rect 8822 10310 8834 10362
rect 8886 10310 8898 10362
rect 8950 10310 8962 10362
rect 9014 10310 9026 10362
rect 9078 10310 11898 10362
rect 11950 10310 11962 10362
rect 12014 10310 12026 10362
rect 12078 10310 12090 10362
rect 12142 10310 12154 10362
rect 12206 10310 13616 10362
rect 1104 10288 13616 10310
rect 6270 10248 6276 10260
rect 4264 10220 6276 10248
rect 4065 10047 4123 10053
rect 4065 10013 4077 10047
rect 4111 10044 4123 10047
rect 4264 10044 4292 10220
rect 6270 10208 6276 10220
rect 6328 10208 6334 10260
rect 6914 10208 6920 10260
rect 6972 10248 6978 10260
rect 7650 10248 7656 10260
rect 6972 10220 7656 10248
rect 6972 10208 6978 10220
rect 7650 10208 7656 10220
rect 7708 10208 7714 10260
rect 4430 10072 4436 10124
rect 4488 10112 4494 10124
rect 8110 10112 8116 10124
rect 4488 10084 8116 10112
rect 4488 10072 4494 10084
rect 4540 10053 4568 10084
rect 8110 10072 8116 10084
rect 8168 10072 8174 10124
rect 9766 10112 9772 10124
rect 9727 10084 9772 10112
rect 9766 10072 9772 10084
rect 9824 10072 9830 10124
rect 10410 10072 10416 10124
rect 10468 10112 10474 10124
rect 11241 10115 11299 10121
rect 11241 10112 11253 10115
rect 10468 10084 11253 10112
rect 10468 10072 10474 10084
rect 11241 10081 11253 10084
rect 11287 10112 11299 10115
rect 12618 10112 12624 10124
rect 11287 10084 12624 10112
rect 11287 10081 11299 10084
rect 11241 10075 11299 10081
rect 12618 10072 12624 10084
rect 12676 10072 12682 10124
rect 12713 10115 12771 10121
rect 12713 10081 12725 10115
rect 12759 10112 12771 10115
rect 12802 10112 12808 10124
rect 12759 10084 12808 10112
rect 12759 10081 12771 10084
rect 12713 10075 12771 10081
rect 12802 10072 12808 10084
rect 12860 10072 12866 10124
rect 4111 10016 4292 10044
rect 4341 10047 4399 10053
rect 4111 10013 4123 10016
rect 4065 10007 4123 10013
rect 4341 10013 4353 10047
rect 4387 10013 4399 10047
rect 4341 10007 4399 10013
rect 4525 10047 4583 10053
rect 4525 10013 4537 10047
rect 4571 10013 4583 10047
rect 4525 10007 4583 10013
rect 4356 9976 4384 10007
rect 4614 10004 4620 10056
rect 4672 10044 4678 10056
rect 4982 10044 4988 10056
rect 4672 10016 4988 10044
rect 4672 10004 4678 10016
rect 4982 10004 4988 10016
rect 5040 10004 5046 10056
rect 5905 10047 5963 10053
rect 5905 10013 5917 10047
rect 5951 10013 5963 10047
rect 9490 10044 9496 10056
rect 9451 10016 9496 10044
rect 5905 10007 5963 10013
rect 5920 9976 5948 10007
rect 9490 10004 9496 10016
rect 9548 10004 9554 10056
rect 12434 10044 12440 10056
rect 12395 10016 12440 10044
rect 12434 10004 12440 10016
rect 12492 10004 12498 10056
rect 6181 9979 6239 9985
rect 4356 9948 4568 9976
rect 5920 9948 6040 9976
rect 4540 9920 4568 9948
rect 3050 9868 3056 9920
rect 3108 9908 3114 9920
rect 3881 9911 3939 9917
rect 3881 9908 3893 9911
rect 3108 9880 3893 9908
rect 3108 9868 3114 9880
rect 3881 9877 3893 9880
rect 3927 9877 3939 9911
rect 3881 9871 3939 9877
rect 4522 9868 4528 9920
rect 4580 9868 4586 9920
rect 5169 9911 5227 9917
rect 5169 9877 5181 9911
rect 5215 9908 5227 9911
rect 6012 9908 6040 9948
rect 6181 9945 6193 9979
rect 6227 9976 6239 9979
rect 6270 9976 6276 9988
rect 6227 9948 6276 9976
rect 6227 9945 6239 9948
rect 6181 9939 6239 9945
rect 6270 9936 6276 9948
rect 6328 9936 6334 9988
rect 6914 9936 6920 9988
rect 6972 9936 6978 9988
rect 12710 9976 12716 9988
rect 10994 9948 12716 9976
rect 12710 9936 12716 9948
rect 12768 9936 12774 9988
rect 6546 9908 6552 9920
rect 5215 9880 6552 9908
rect 5215 9877 5227 9880
rect 5169 9871 5227 9877
rect 6546 9868 6552 9880
rect 6604 9868 6610 9920
rect 12069 9911 12127 9917
rect 12069 9877 12081 9911
rect 12115 9908 12127 9911
rect 12158 9908 12164 9920
rect 12115 9880 12164 9908
rect 12115 9877 12127 9880
rect 12069 9871 12127 9877
rect 12158 9868 12164 9880
rect 12216 9868 12222 9920
rect 12526 9868 12532 9920
rect 12584 9908 12590 9920
rect 12584 9880 12629 9908
rect 12584 9868 12590 9880
rect 1104 9818 13616 9840
rect 1104 9766 4078 9818
rect 4130 9766 4142 9818
rect 4194 9766 4206 9818
rect 4258 9766 4270 9818
rect 4322 9766 4334 9818
rect 4386 9766 7206 9818
rect 7258 9766 7270 9818
rect 7322 9766 7334 9818
rect 7386 9766 7398 9818
rect 7450 9766 7462 9818
rect 7514 9766 10334 9818
rect 10386 9766 10398 9818
rect 10450 9766 10462 9818
rect 10514 9766 10526 9818
rect 10578 9766 10590 9818
rect 10642 9766 13616 9818
rect 1104 9744 13616 9766
rect 4249 9639 4307 9645
rect 4249 9605 4261 9639
rect 4295 9636 4307 9639
rect 4522 9636 4528 9648
rect 4295 9608 4528 9636
rect 4295 9605 4307 9608
rect 4249 9599 4307 9605
rect 4522 9596 4528 9608
rect 4580 9596 4586 9648
rect 6733 9639 6791 9645
rect 6733 9636 6745 9639
rect 5474 9622 6745 9636
rect 5460 9608 6745 9622
rect 2866 9528 2872 9580
rect 2924 9528 2930 9580
rect 1394 9460 1400 9512
rect 1452 9500 1458 9512
rect 1489 9503 1547 9509
rect 1489 9500 1501 9503
rect 1452 9472 1501 9500
rect 1452 9460 1458 9472
rect 1489 9469 1501 9472
rect 1535 9469 1547 9503
rect 1762 9500 1768 9512
rect 1723 9472 1768 9500
rect 1489 9463 1547 9469
rect 1762 9460 1768 9472
rect 1820 9460 1826 9512
rect 2884 9432 2912 9528
rect 3234 9500 3240 9512
rect 3195 9472 3240 9500
rect 3234 9460 3240 9472
rect 3292 9460 3298 9512
rect 3970 9500 3976 9512
rect 3931 9472 3976 9500
rect 3970 9460 3976 9472
rect 4028 9460 4034 9512
rect 5460 9500 5488 9608
rect 6733 9605 6745 9608
rect 6779 9605 6791 9639
rect 6733 9599 6791 9605
rect 6914 9528 6920 9580
rect 6972 9568 6978 9580
rect 9217 9571 9275 9577
rect 6972 9540 7017 9568
rect 6972 9528 6978 9540
rect 9217 9537 9229 9571
rect 9263 9568 9275 9571
rect 9306 9568 9312 9580
rect 9263 9540 9312 9568
rect 9263 9537 9275 9540
rect 9217 9531 9275 9537
rect 9306 9528 9312 9540
rect 9364 9528 9370 9580
rect 12158 9568 12164 9580
rect 12119 9540 12164 9568
rect 12158 9528 12164 9540
rect 12216 9528 12222 9580
rect 9030 9500 9036 9512
rect 4080 9472 5488 9500
rect 8991 9472 9036 9500
rect 4080 9432 4108 9472
rect 9030 9460 9036 9472
rect 9088 9460 9094 9512
rect 9125 9503 9183 9509
rect 9125 9469 9137 9503
rect 9171 9469 9183 9503
rect 9125 9463 9183 9469
rect 2884 9404 4108 9432
rect 5350 9392 5356 9444
rect 5408 9432 5414 9444
rect 9140 9432 9168 9463
rect 5408 9404 9168 9432
rect 9585 9435 9643 9441
rect 5408 9392 5414 9404
rect 9585 9401 9597 9435
rect 9631 9432 9643 9435
rect 9950 9432 9956 9444
rect 9631 9404 9956 9432
rect 9631 9401 9643 9404
rect 9585 9395 9643 9401
rect 9950 9392 9956 9404
rect 10008 9392 10014 9444
rect 5258 9324 5264 9376
rect 5316 9364 5322 9376
rect 5721 9367 5779 9373
rect 5721 9364 5733 9367
rect 5316 9336 5733 9364
rect 5316 9324 5322 9336
rect 5721 9333 5733 9336
rect 5767 9333 5779 9367
rect 5721 9327 5779 9333
rect 11422 9324 11428 9376
rect 11480 9364 11486 9376
rect 11977 9367 12035 9373
rect 11977 9364 11989 9367
rect 11480 9336 11989 9364
rect 11480 9324 11486 9336
rect 11977 9333 11989 9336
rect 12023 9333 12035 9367
rect 11977 9327 12035 9333
rect 1104 9274 13616 9296
rect 1104 9222 2514 9274
rect 2566 9222 2578 9274
rect 2630 9222 2642 9274
rect 2694 9222 2706 9274
rect 2758 9222 2770 9274
rect 2822 9222 5642 9274
rect 5694 9222 5706 9274
rect 5758 9222 5770 9274
rect 5822 9222 5834 9274
rect 5886 9222 5898 9274
rect 5950 9222 8770 9274
rect 8822 9222 8834 9274
rect 8886 9222 8898 9274
rect 8950 9222 8962 9274
rect 9014 9222 9026 9274
rect 9078 9222 11898 9274
rect 11950 9222 11962 9274
rect 12014 9222 12026 9274
rect 12078 9222 12090 9274
rect 12142 9222 12154 9274
rect 12206 9222 13616 9274
rect 1104 9200 13616 9222
rect 1762 9120 1768 9172
rect 1820 9160 1826 9172
rect 2593 9163 2651 9169
rect 2593 9160 2605 9163
rect 1820 9132 2605 9160
rect 1820 9120 1826 9132
rect 2593 9129 2605 9132
rect 2639 9129 2651 9163
rect 6270 9160 6276 9172
rect 2593 9123 2651 9129
rect 5092 9132 6276 9160
rect 3789 9095 3847 9101
rect 3789 9061 3801 9095
rect 3835 9061 3847 9095
rect 3789 9055 3847 9061
rect 3804 9024 3832 9055
rect 2792 8996 3832 9024
rect 4433 9027 4491 9033
rect 2792 8965 2820 8996
rect 4433 8993 4445 9027
rect 4479 9024 4491 9027
rect 5092 9024 5120 9132
rect 6270 9120 6276 9132
rect 6328 9160 6334 9172
rect 6733 9163 6791 9169
rect 6733 9160 6745 9163
rect 6328 9132 6745 9160
rect 6328 9120 6334 9132
rect 6733 9129 6745 9132
rect 6779 9129 6791 9163
rect 6733 9123 6791 9129
rect 12434 9120 12440 9172
rect 12492 9160 12498 9172
rect 12897 9163 12955 9169
rect 12897 9160 12909 9163
rect 12492 9132 12909 9160
rect 12492 9120 12498 9132
rect 12897 9129 12909 9132
rect 12943 9129 12955 9163
rect 12897 9123 12955 9129
rect 5258 9024 5264 9036
rect 4479 8996 5120 9024
rect 5219 8996 5264 9024
rect 4479 8993 4491 8996
rect 4433 8987 4491 8993
rect 5258 8984 5264 8996
rect 5316 8984 5322 9036
rect 11422 9024 11428 9036
rect 11383 8996 11428 9024
rect 11422 8984 11428 8996
rect 11480 8984 11486 9036
rect 2777 8959 2835 8965
rect 2777 8925 2789 8959
rect 2823 8925 2835 8959
rect 3050 8956 3056 8968
rect 3011 8928 3056 8956
rect 2777 8919 2835 8925
rect 3050 8916 3056 8928
rect 3108 8916 3114 8968
rect 3234 8956 3240 8968
rect 3195 8928 3240 8956
rect 3234 8916 3240 8928
rect 3292 8916 3298 8968
rect 4982 8956 4988 8968
rect 4943 8928 4988 8956
rect 4982 8916 4988 8928
rect 5040 8916 5046 8968
rect 9490 8916 9496 8968
rect 9548 8956 9554 8968
rect 10226 8956 10232 8968
rect 9548 8928 10232 8956
rect 9548 8916 9554 8928
rect 10226 8916 10232 8928
rect 10284 8956 10290 8968
rect 11149 8959 11207 8965
rect 11149 8956 11161 8959
rect 10284 8928 11161 8956
rect 10284 8916 10290 8928
rect 11149 8925 11161 8928
rect 11195 8925 11207 8959
rect 11149 8919 11207 8925
rect 4157 8891 4215 8897
rect 4157 8857 4169 8891
rect 4203 8888 4215 8891
rect 4614 8888 4620 8900
rect 4203 8860 4620 8888
rect 4203 8857 4215 8860
rect 4157 8851 4215 8857
rect 4614 8848 4620 8860
rect 4672 8848 4678 8900
rect 6914 8888 6920 8900
rect 6486 8860 6920 8888
rect 6914 8848 6920 8860
rect 6972 8888 6978 8900
rect 7558 8888 7564 8900
rect 6972 8860 7564 8888
rect 6972 8848 6978 8860
rect 7558 8848 7564 8860
rect 7616 8848 7622 8900
rect 4249 8823 4307 8829
rect 4249 8789 4261 8823
rect 4295 8820 4307 8823
rect 4706 8820 4712 8832
rect 4295 8792 4712 8820
rect 4295 8789 4307 8792
rect 4249 8783 4307 8789
rect 4706 8780 4712 8792
rect 4764 8820 4770 8832
rect 5350 8820 5356 8832
rect 4764 8792 5356 8820
rect 4764 8780 4770 8792
rect 5350 8780 5356 8792
rect 5408 8780 5414 8832
rect 11164 8820 11192 8919
rect 12710 8888 12716 8900
rect 12650 8860 12716 8888
rect 12710 8848 12716 8860
rect 12768 8848 12774 8900
rect 12894 8820 12900 8832
rect 11164 8792 12900 8820
rect 12894 8780 12900 8792
rect 12952 8780 12958 8832
rect 1104 8730 13616 8752
rect 1104 8678 4078 8730
rect 4130 8678 4142 8730
rect 4194 8678 4206 8730
rect 4258 8678 4270 8730
rect 4322 8678 4334 8730
rect 4386 8678 7206 8730
rect 7258 8678 7270 8730
rect 7322 8678 7334 8730
rect 7386 8678 7398 8730
rect 7450 8678 7462 8730
rect 7514 8678 10334 8730
rect 10386 8678 10398 8730
rect 10450 8678 10462 8730
rect 10514 8678 10526 8730
rect 10578 8678 10590 8730
rect 10642 8678 13616 8730
rect 1104 8656 13616 8678
rect 4157 8619 4215 8625
rect 4157 8585 4169 8619
rect 4203 8616 4215 8619
rect 4982 8616 4988 8628
rect 4203 8588 4988 8616
rect 4203 8585 4215 8588
rect 4157 8579 4215 8585
rect 4982 8576 4988 8588
rect 5040 8576 5046 8628
rect 9490 8576 9496 8628
rect 9548 8616 9554 8628
rect 9585 8619 9643 8625
rect 9585 8616 9597 8619
rect 9548 8588 9597 8616
rect 9548 8576 9554 8588
rect 9585 8585 9597 8588
rect 9631 8585 9643 8619
rect 12802 8616 12808 8628
rect 12763 8588 12808 8616
rect 9585 8579 9643 8585
rect 12802 8576 12808 8588
rect 12860 8576 12866 8628
rect 3970 8480 3976 8492
rect 3931 8452 3976 8480
rect 3970 8440 3976 8452
rect 4028 8440 4034 8492
rect 9122 8440 9128 8492
rect 9180 8480 9186 8492
rect 9401 8483 9459 8489
rect 9401 8480 9413 8483
rect 9180 8452 9413 8480
rect 9180 8440 9186 8452
rect 9401 8449 9413 8452
rect 9447 8449 9459 8483
rect 12618 8480 12624 8492
rect 12579 8452 12624 8480
rect 9401 8443 9459 8449
rect 12618 8440 12624 8452
rect 12676 8440 12682 8492
rect 1104 8186 13616 8208
rect 1104 8134 2514 8186
rect 2566 8134 2578 8186
rect 2630 8134 2642 8186
rect 2694 8134 2706 8186
rect 2758 8134 2770 8186
rect 2822 8134 5642 8186
rect 5694 8134 5706 8186
rect 5758 8134 5770 8186
rect 5822 8134 5834 8186
rect 5886 8134 5898 8186
rect 5950 8134 8770 8186
rect 8822 8134 8834 8186
rect 8886 8134 8898 8186
rect 8950 8134 8962 8186
rect 9014 8134 9026 8186
rect 9078 8134 11898 8186
rect 11950 8134 11962 8186
rect 12014 8134 12026 8186
rect 12078 8134 12090 8186
rect 12142 8134 12154 8186
rect 12206 8134 13616 8186
rect 1104 8112 13616 8134
rect 11149 8075 11207 8081
rect 11149 8072 11161 8075
rect 7944 8044 11161 8072
rect 7006 7896 7012 7948
rect 7064 7936 7070 7948
rect 7064 7908 7328 7936
rect 7064 7896 7070 7908
rect 1673 7871 1731 7877
rect 1673 7837 1685 7871
rect 1719 7868 1731 7871
rect 2038 7868 2044 7880
rect 1719 7840 2044 7868
rect 1719 7837 1731 7840
rect 1673 7831 1731 7837
rect 2038 7828 2044 7840
rect 2096 7828 2102 7880
rect 2314 7868 2320 7880
rect 2275 7840 2320 7868
rect 2314 7828 2320 7840
rect 2372 7828 2378 7880
rect 3789 7871 3847 7877
rect 3789 7837 3801 7871
rect 3835 7868 3847 7871
rect 3970 7868 3976 7880
rect 3835 7840 3976 7868
rect 3835 7837 3847 7840
rect 3789 7831 3847 7837
rect 3970 7828 3976 7840
rect 4028 7828 4034 7880
rect 6825 7871 6883 7877
rect 6825 7837 6837 7871
rect 6871 7868 6883 7871
rect 6914 7868 6920 7880
rect 6871 7840 6920 7868
rect 6871 7837 6883 7840
rect 6825 7831 6883 7837
rect 6914 7828 6920 7840
rect 6972 7828 6978 7880
rect 7300 7877 7328 7908
rect 7101 7871 7159 7877
rect 7101 7837 7113 7871
rect 7147 7837 7159 7871
rect 7101 7831 7159 7837
rect 7285 7871 7343 7877
rect 7285 7837 7297 7871
rect 7331 7837 7343 7871
rect 7285 7831 7343 7837
rect 7116 7800 7144 7831
rect 7650 7828 7656 7880
rect 7708 7868 7714 7880
rect 7944 7877 7972 8044
rect 11149 8041 11161 8044
rect 11195 8041 11207 8075
rect 11149 8035 11207 8041
rect 9217 7939 9275 7945
rect 9217 7936 9229 7939
rect 8404 7908 9229 7936
rect 7929 7871 7987 7877
rect 7929 7868 7941 7871
rect 7708 7840 7941 7868
rect 7708 7828 7714 7840
rect 7929 7837 7941 7840
rect 7975 7837 7987 7871
rect 7929 7831 7987 7837
rect 8205 7871 8263 7877
rect 8205 7837 8217 7871
rect 8251 7837 8263 7871
rect 8205 7831 8263 7837
rect 7745 7803 7803 7809
rect 7745 7800 7757 7803
rect 7116 7772 7757 7800
rect 7745 7769 7757 7772
rect 7791 7769 7803 7803
rect 8220 7800 8248 7831
rect 8294 7828 8300 7880
rect 8352 7868 8358 7880
rect 8404 7877 8432 7908
rect 9217 7905 9229 7908
rect 9263 7905 9275 7939
rect 12894 7936 12900 7948
rect 12855 7908 12900 7936
rect 9217 7899 9275 7905
rect 12894 7896 12900 7908
rect 12952 7896 12958 7948
rect 8389 7871 8447 7877
rect 8389 7868 8401 7871
rect 8352 7840 8401 7868
rect 8352 7828 8358 7840
rect 8389 7837 8401 7840
rect 8435 7837 8447 7871
rect 8938 7868 8944 7880
rect 8899 7840 8944 7868
rect 8389 7831 8447 7837
rect 8938 7828 8944 7840
rect 8996 7828 9002 7880
rect 9490 7800 9496 7812
rect 8220 7772 9496 7800
rect 7745 7763 7803 7769
rect 9490 7760 9496 7772
rect 9548 7760 9554 7812
rect 9600 7772 9706 7800
rect 12190 7772 12296 7800
rect 9600 7744 9628 7772
rect 1486 7732 1492 7744
rect 1447 7704 1492 7732
rect 1486 7692 1492 7704
rect 1544 7692 1550 7744
rect 1670 7692 1676 7744
rect 1728 7732 1734 7744
rect 2133 7735 2191 7741
rect 2133 7732 2145 7735
rect 1728 7704 2145 7732
rect 1728 7692 1734 7704
rect 2133 7701 2145 7704
rect 2179 7701 2191 7735
rect 2133 7695 2191 7701
rect 3973 7735 4031 7741
rect 3973 7701 3985 7735
rect 4019 7732 4031 7735
rect 4430 7732 4436 7744
rect 4019 7704 4436 7732
rect 4019 7701 4031 7704
rect 3973 7695 4031 7701
rect 4430 7692 4436 7704
rect 4488 7692 4494 7744
rect 6638 7732 6644 7744
rect 6599 7704 6644 7732
rect 6638 7692 6644 7704
rect 6696 7692 6702 7744
rect 7098 7692 7104 7744
rect 7156 7732 7162 7744
rect 9582 7732 9588 7744
rect 7156 7704 9588 7732
rect 7156 7692 7162 7704
rect 9582 7692 9588 7704
rect 9640 7692 9646 7744
rect 10686 7732 10692 7744
rect 10647 7704 10692 7732
rect 10686 7692 10692 7704
rect 10744 7692 10750 7744
rect 12268 7732 12296 7772
rect 12342 7760 12348 7812
rect 12400 7800 12406 7812
rect 12621 7803 12679 7809
rect 12621 7800 12633 7803
rect 12400 7772 12633 7800
rect 12400 7760 12406 7772
rect 12621 7769 12633 7772
rect 12667 7769 12679 7803
rect 12621 7763 12679 7769
rect 12802 7732 12808 7744
rect 12268 7704 12808 7732
rect 12802 7692 12808 7704
rect 12860 7692 12866 7744
rect 1104 7642 13616 7664
rect 1104 7590 4078 7642
rect 4130 7590 4142 7642
rect 4194 7590 4206 7642
rect 4258 7590 4270 7642
rect 4322 7590 4334 7642
rect 4386 7590 7206 7642
rect 7258 7590 7270 7642
rect 7322 7590 7334 7642
rect 7386 7590 7398 7642
rect 7450 7590 7462 7642
rect 7514 7590 10334 7642
rect 10386 7590 10398 7642
rect 10450 7590 10462 7642
rect 10514 7590 10526 7642
rect 10578 7590 10590 7642
rect 10642 7590 13616 7642
rect 1104 7568 13616 7590
rect 2038 7488 2044 7540
rect 2096 7528 2102 7540
rect 3145 7531 3203 7537
rect 3145 7528 3157 7531
rect 2096 7500 3157 7528
rect 2096 7488 2102 7500
rect 3145 7497 3157 7500
rect 3191 7497 3203 7531
rect 3145 7491 3203 7497
rect 7558 7488 7564 7540
rect 7616 7528 7622 7540
rect 8573 7531 8631 7537
rect 8573 7528 8585 7531
rect 7616 7500 8585 7528
rect 7616 7488 7622 7500
rect 8573 7497 8585 7500
rect 8619 7497 8631 7531
rect 8573 7491 8631 7497
rect 9490 7488 9496 7540
rect 9548 7528 9554 7540
rect 10962 7528 10968 7540
rect 9548 7500 10968 7528
rect 9548 7488 9554 7500
rect 10962 7488 10968 7500
rect 11020 7488 11026 7540
rect 12710 7528 12716 7540
rect 12671 7500 12716 7528
rect 12710 7488 12716 7500
rect 12768 7488 12774 7540
rect 1670 7460 1676 7472
rect 1631 7432 1676 7460
rect 1670 7420 1676 7432
rect 1728 7420 1734 7472
rect 3878 7460 3884 7472
rect 2898 7432 3884 7460
rect 3878 7420 3884 7432
rect 3936 7420 3942 7472
rect 6638 7460 6644 7472
rect 6599 7432 6644 7460
rect 6638 7420 6644 7432
rect 6696 7420 6702 7472
rect 7098 7420 7104 7472
rect 7156 7420 7162 7472
rect 9582 7420 9588 7472
rect 9640 7460 9646 7472
rect 9640 7432 9982 7460
rect 9640 7420 9646 7432
rect 3602 7392 3608 7404
rect 3515 7364 3608 7392
rect 3602 7352 3608 7364
rect 3660 7392 3666 7404
rect 3970 7392 3976 7404
rect 3660 7364 3976 7392
rect 3660 7352 3666 7364
rect 3970 7352 3976 7364
rect 4028 7352 4034 7404
rect 4430 7392 4436 7404
rect 4391 7364 4436 7392
rect 4430 7352 4436 7364
rect 4488 7392 4494 7404
rect 4890 7392 4896 7404
rect 4488 7364 4896 7392
rect 4488 7352 4494 7364
rect 4890 7352 4896 7364
rect 4948 7352 4954 7404
rect 8294 7352 8300 7404
rect 8352 7392 8358 7404
rect 8757 7395 8815 7401
rect 8757 7392 8769 7395
rect 8352 7364 8769 7392
rect 8352 7352 8358 7364
rect 8757 7361 8769 7364
rect 8803 7361 8815 7395
rect 8757 7355 8815 7361
rect 12069 7395 12127 7401
rect 12069 7361 12081 7395
rect 12115 7392 12127 7395
rect 12802 7392 12808 7404
rect 12115 7364 12808 7392
rect 12115 7361 12127 7364
rect 12069 7355 12127 7361
rect 12802 7352 12808 7364
rect 12860 7352 12866 7404
rect 1394 7324 1400 7336
rect 1307 7296 1400 7324
rect 1394 7284 1400 7296
rect 1452 7284 1458 7336
rect 6365 7327 6423 7333
rect 6365 7293 6377 7327
rect 6411 7324 6423 7327
rect 8938 7324 8944 7336
rect 6411 7296 8944 7324
rect 6411 7293 6423 7296
rect 6365 7287 6423 7293
rect 1412 7188 1440 7284
rect 3789 7259 3847 7265
rect 3789 7225 3801 7259
rect 3835 7256 3847 7259
rect 6380 7256 6408 7287
rect 8938 7284 8944 7296
rect 8996 7324 9002 7336
rect 9217 7327 9275 7333
rect 9217 7324 9229 7327
rect 8996 7296 9229 7324
rect 8996 7284 9002 7296
rect 9217 7293 9229 7296
rect 9263 7293 9275 7327
rect 9217 7287 9275 7293
rect 9493 7327 9551 7333
rect 9493 7293 9505 7327
rect 9539 7324 9551 7327
rect 9858 7324 9864 7336
rect 9539 7296 9864 7324
rect 9539 7293 9551 7296
rect 9493 7287 9551 7293
rect 9858 7284 9864 7296
rect 9916 7324 9922 7336
rect 10686 7324 10692 7336
rect 9916 7296 10692 7324
rect 9916 7284 9922 7296
rect 10686 7284 10692 7296
rect 10744 7284 10750 7336
rect 3835 7228 6408 7256
rect 3835 7225 3847 7228
rect 3789 7219 3847 7225
rect 4249 7191 4307 7197
rect 4249 7188 4261 7191
rect 1412 7160 4261 7188
rect 4249 7157 4261 7160
rect 4295 7157 4307 7191
rect 4249 7151 4307 7157
rect 7006 7148 7012 7200
rect 7064 7188 7070 7200
rect 8113 7191 8171 7197
rect 8113 7188 8125 7191
rect 7064 7160 8125 7188
rect 7064 7148 7070 7160
rect 8113 7157 8125 7160
rect 8159 7157 8171 7191
rect 8113 7151 8171 7157
rect 9582 7148 9588 7200
rect 9640 7188 9646 7200
rect 11977 7191 12035 7197
rect 11977 7188 11989 7191
rect 9640 7160 11989 7188
rect 9640 7148 9646 7160
rect 11977 7157 11989 7160
rect 12023 7157 12035 7191
rect 11977 7151 12035 7157
rect 1104 7098 13616 7120
rect 1104 7046 2514 7098
rect 2566 7046 2578 7098
rect 2630 7046 2642 7098
rect 2694 7046 2706 7098
rect 2758 7046 2770 7098
rect 2822 7046 5642 7098
rect 5694 7046 5706 7098
rect 5758 7046 5770 7098
rect 5822 7046 5834 7098
rect 5886 7046 5898 7098
rect 5950 7046 8770 7098
rect 8822 7046 8834 7098
rect 8886 7046 8898 7098
rect 8950 7046 8962 7098
rect 9014 7046 9026 7098
rect 9078 7046 11898 7098
rect 11950 7046 11962 7098
rect 12014 7046 12026 7098
rect 12078 7046 12090 7098
rect 12142 7046 12154 7098
rect 12206 7046 13616 7098
rect 1104 7024 13616 7046
rect 2314 6984 2320 6996
rect 2275 6956 2320 6984
rect 2314 6944 2320 6956
rect 2372 6944 2378 6996
rect 3970 6944 3976 6996
rect 4028 6984 4034 6996
rect 4230 6987 4288 6993
rect 4230 6984 4242 6987
rect 4028 6956 4242 6984
rect 4028 6944 4034 6956
rect 4230 6953 4242 6956
rect 4276 6953 4288 6987
rect 4230 6947 4288 6953
rect 6914 6944 6920 6996
rect 6972 6984 6978 6996
rect 6972 6956 7017 6984
rect 6972 6944 6978 6956
rect 9858 6916 9864 6928
rect 9508 6888 9864 6916
rect 2406 6808 2412 6860
rect 2464 6848 2470 6860
rect 2869 6851 2927 6857
rect 2869 6848 2881 6851
rect 2464 6820 2881 6848
rect 2464 6808 2470 6820
rect 2869 6817 2881 6820
rect 2915 6817 2927 6851
rect 2869 6811 2927 6817
rect 3973 6851 4031 6857
rect 3973 6817 3985 6851
rect 4019 6848 4031 6851
rect 4890 6848 4896 6860
rect 4019 6820 4896 6848
rect 4019 6817 4031 6820
rect 3973 6811 4031 6817
rect 4890 6808 4896 6820
rect 4948 6808 4954 6860
rect 5258 6808 5264 6860
rect 5316 6848 5322 6860
rect 7558 6848 7564 6860
rect 5316 6820 6914 6848
rect 7519 6820 7564 6848
rect 5316 6808 5322 6820
rect 2038 6740 2044 6792
rect 2096 6780 2102 6792
rect 2685 6783 2743 6789
rect 2685 6780 2697 6783
rect 2096 6752 2697 6780
rect 2096 6740 2102 6752
rect 2685 6749 2697 6752
rect 2731 6749 2743 6783
rect 6886 6780 6914 6820
rect 7558 6808 7564 6820
rect 7616 6808 7622 6860
rect 9217 6851 9275 6857
rect 9217 6817 9229 6851
rect 9263 6848 9275 6851
rect 9508 6848 9536 6888
rect 9858 6876 9864 6888
rect 9916 6876 9922 6928
rect 9263 6820 9536 6848
rect 9263 6817 9275 6820
rect 9217 6811 9275 6817
rect 10226 6808 10232 6860
rect 10284 6848 10290 6860
rect 10505 6851 10563 6857
rect 10505 6848 10517 6851
rect 10284 6820 10517 6848
rect 10284 6808 10290 6820
rect 10505 6817 10517 6820
rect 10551 6817 10563 6851
rect 10505 6811 10563 6817
rect 10781 6851 10839 6857
rect 10781 6817 10793 6851
rect 10827 6848 10839 6851
rect 10870 6848 10876 6860
rect 10827 6820 10876 6848
rect 10827 6817 10839 6820
rect 10781 6811 10839 6817
rect 10870 6808 10876 6820
rect 10928 6808 10934 6860
rect 12253 6851 12311 6857
rect 12253 6817 12265 6851
rect 12299 6848 12311 6851
rect 12342 6848 12348 6860
rect 12299 6820 12348 6848
rect 12299 6817 12311 6820
rect 12253 6811 12311 6817
rect 12342 6808 12348 6820
rect 12400 6808 12406 6860
rect 7285 6783 7343 6789
rect 7285 6780 7297 6783
rect 6886 6752 7297 6780
rect 2685 6743 2743 6749
rect 7285 6749 7297 6752
rect 7331 6780 7343 6783
rect 8570 6780 8576 6792
rect 7331 6752 8576 6780
rect 7331 6749 7343 6752
rect 7285 6743 7343 6749
rect 8570 6740 8576 6752
rect 8628 6780 8634 6792
rect 9306 6780 9312 6792
rect 8628 6752 9312 6780
rect 8628 6740 8634 6752
rect 9306 6740 9312 6752
rect 9364 6780 9370 6792
rect 9493 6783 9551 6789
rect 9493 6780 9505 6783
rect 9364 6752 9505 6780
rect 9364 6740 9370 6752
rect 9493 6749 9505 6752
rect 9539 6749 9551 6783
rect 9493 6743 9551 6749
rect 8294 6712 8300 6724
rect 5474 6684 8300 6712
rect 2777 6647 2835 6653
rect 2777 6613 2789 6647
rect 2823 6644 2835 6647
rect 3510 6644 3516 6656
rect 2823 6616 3516 6644
rect 2823 6613 2835 6616
rect 2777 6607 2835 6613
rect 3510 6604 3516 6616
rect 3568 6604 3574 6656
rect 3878 6604 3884 6656
rect 3936 6644 3942 6656
rect 5552 6644 5580 6684
rect 8294 6672 8300 6684
rect 8352 6672 8358 6724
rect 12802 6712 12808 6724
rect 12006 6684 12808 6712
rect 12802 6672 12808 6684
rect 12860 6672 12866 6724
rect 5718 6644 5724 6656
rect 3936 6616 5580 6644
rect 5679 6616 5724 6644
rect 3936 6604 3942 6616
rect 5718 6604 5724 6616
rect 5776 6604 5782 6656
rect 7377 6647 7435 6653
rect 7377 6613 7389 6647
rect 7423 6644 7435 6647
rect 7650 6644 7656 6656
rect 7423 6616 7656 6644
rect 7423 6613 7435 6616
rect 7377 6607 7435 6613
rect 7650 6604 7656 6616
rect 7708 6604 7714 6656
rect 1104 6554 13616 6576
rect 1104 6502 4078 6554
rect 4130 6502 4142 6554
rect 4194 6502 4206 6554
rect 4258 6502 4270 6554
rect 4322 6502 4334 6554
rect 4386 6502 7206 6554
rect 7258 6502 7270 6554
rect 7322 6502 7334 6554
rect 7386 6502 7398 6554
rect 7450 6502 7462 6554
rect 7514 6502 10334 6554
rect 10386 6502 10398 6554
rect 10450 6502 10462 6554
rect 10514 6502 10526 6554
rect 10578 6502 10590 6554
rect 10642 6502 13616 6554
rect 1104 6480 13616 6502
rect 3145 6443 3203 6449
rect 3145 6409 3157 6443
rect 3191 6440 3203 6443
rect 4522 6440 4528 6452
rect 3191 6412 4528 6440
rect 3191 6409 3203 6412
rect 3145 6403 3203 6409
rect 4522 6400 4528 6412
rect 4580 6400 4586 6452
rect 4614 6400 4620 6452
rect 4672 6440 4678 6452
rect 5258 6440 5264 6452
rect 4672 6412 5264 6440
rect 4672 6400 4678 6412
rect 5258 6400 5264 6412
rect 5316 6400 5322 6452
rect 5718 6400 5724 6452
rect 5776 6440 5782 6452
rect 7193 6443 7251 6449
rect 5776 6412 7052 6440
rect 5776 6400 5782 6412
rect 3878 6332 3884 6384
rect 3936 6332 3942 6384
rect 4706 6332 4712 6384
rect 4764 6372 4770 6384
rect 4764 6344 6914 6372
rect 4764 6332 4770 6344
rect 4890 6264 4896 6316
rect 4948 6304 4954 6316
rect 4948 6276 4993 6304
rect 4948 6264 4954 6276
rect 4614 6236 4620 6248
rect 4575 6208 4620 6236
rect 4614 6196 4620 6208
rect 4672 6196 4678 6248
rect 5718 6128 5724 6180
rect 5776 6128 5782 6180
rect 6886 6168 6914 6344
rect 7024 6236 7052 6412
rect 7193 6409 7205 6443
rect 7239 6440 7251 6443
rect 8294 6440 8300 6452
rect 7239 6412 8300 6440
rect 7239 6409 7251 6412
rect 7193 6403 7251 6409
rect 8294 6400 8300 6412
rect 8352 6400 8358 6452
rect 7098 6332 7104 6384
rect 7156 6372 7162 6384
rect 7285 6375 7343 6381
rect 7285 6372 7297 6375
rect 7156 6344 7297 6372
rect 7156 6332 7162 6344
rect 7285 6341 7297 6344
rect 7331 6341 7343 6375
rect 7285 6335 7343 6341
rect 12986 6236 12992 6248
rect 7024 6208 12992 6236
rect 12986 6196 12992 6208
rect 13044 6196 13050 6248
rect 7650 6168 7656 6180
rect 6886 6140 7656 6168
rect 7650 6128 7656 6140
rect 7708 6128 7714 6180
rect 3510 6060 3516 6112
rect 3568 6100 3574 6112
rect 5534 6100 5540 6112
rect 3568 6072 5540 6100
rect 3568 6060 3574 6072
rect 5534 6060 5540 6072
rect 5592 6100 5598 6112
rect 5736 6100 5764 6128
rect 5592 6072 5764 6100
rect 5592 6060 5598 6072
rect 1104 6010 13616 6032
rect 1104 5958 2514 6010
rect 2566 5958 2578 6010
rect 2630 5958 2642 6010
rect 2694 5958 2706 6010
rect 2758 5958 2770 6010
rect 2822 5958 5642 6010
rect 5694 5958 5706 6010
rect 5758 5958 5770 6010
rect 5822 5958 5834 6010
rect 5886 5958 5898 6010
rect 5950 5958 8770 6010
rect 8822 5958 8834 6010
rect 8886 5958 8898 6010
rect 8950 5958 8962 6010
rect 9014 5958 9026 6010
rect 9078 5958 11898 6010
rect 11950 5958 11962 6010
rect 12014 5958 12026 6010
rect 12078 5958 12090 6010
rect 12142 5958 12154 6010
rect 12206 5958 13616 6010
rect 1104 5936 13616 5958
rect 12802 5828 12808 5840
rect 12763 5800 12808 5828
rect 12802 5788 12808 5800
rect 12860 5788 12866 5840
rect 4525 5763 4583 5769
rect 4525 5729 4537 5763
rect 4571 5760 4583 5763
rect 4614 5760 4620 5772
rect 4571 5732 4620 5760
rect 4571 5729 4583 5732
rect 4525 5723 4583 5729
rect 4614 5720 4620 5732
rect 4672 5760 4678 5772
rect 5166 5760 5172 5772
rect 4672 5732 5172 5760
rect 4672 5720 4678 5732
rect 5166 5720 5172 5732
rect 5224 5720 5230 5772
rect 9674 5760 9680 5772
rect 9635 5732 9680 5760
rect 9674 5720 9680 5732
rect 9732 5720 9738 5772
rect 9858 5652 9864 5704
rect 9916 5692 9922 5704
rect 9953 5695 10011 5701
rect 9953 5692 9965 5695
rect 9916 5664 9965 5692
rect 9916 5652 9922 5664
rect 9953 5661 9965 5664
rect 9999 5661 10011 5695
rect 11057 5695 11115 5701
rect 11057 5692 11069 5695
rect 9953 5655 10011 5661
rect 10336 5664 11069 5692
rect 4249 5627 4307 5633
rect 4249 5593 4261 5627
rect 4295 5624 4307 5627
rect 4522 5624 4528 5636
rect 4295 5596 4528 5624
rect 4295 5593 4307 5596
rect 4249 5587 4307 5593
rect 4522 5584 4528 5596
rect 4580 5584 4586 5636
rect 3878 5556 3884 5568
rect 3839 5528 3884 5556
rect 3878 5516 3884 5528
rect 3936 5516 3942 5568
rect 4341 5559 4399 5565
rect 4341 5525 4353 5559
rect 4387 5556 4399 5559
rect 4430 5556 4436 5568
rect 4387 5528 4436 5556
rect 4387 5525 4399 5528
rect 4341 5519 4399 5525
rect 4430 5516 4436 5528
rect 4488 5556 4494 5568
rect 4706 5556 4712 5568
rect 4488 5528 4712 5556
rect 4488 5516 4494 5528
rect 4706 5516 4712 5528
rect 4764 5516 4770 5568
rect 7650 5516 7656 5568
rect 7708 5556 7714 5568
rect 10336 5565 10364 5664
rect 11057 5661 11069 5664
rect 11103 5661 11115 5695
rect 11330 5692 11336 5704
rect 11291 5664 11336 5692
rect 11057 5655 11115 5661
rect 11330 5652 11336 5664
rect 11388 5652 11394 5704
rect 11517 5695 11575 5701
rect 11517 5661 11529 5695
rect 11563 5692 11575 5695
rect 12526 5692 12532 5704
rect 11563 5664 12532 5692
rect 11563 5661 11575 5664
rect 11517 5655 11575 5661
rect 12526 5652 12532 5664
rect 12584 5692 12590 5704
rect 12802 5692 12808 5704
rect 12584 5664 12808 5692
rect 12584 5652 12590 5664
rect 12802 5652 12808 5664
rect 12860 5652 12866 5704
rect 12618 5624 12624 5636
rect 12579 5596 12624 5624
rect 12618 5584 12624 5596
rect 12676 5584 12682 5636
rect 9861 5559 9919 5565
rect 9861 5556 9873 5559
rect 7708 5528 9873 5556
rect 7708 5516 7714 5528
rect 9861 5525 9873 5528
rect 9907 5525 9919 5559
rect 9861 5519 9919 5525
rect 10321 5559 10379 5565
rect 10321 5525 10333 5559
rect 10367 5525 10379 5559
rect 10321 5519 10379 5525
rect 10873 5559 10931 5565
rect 10873 5525 10885 5559
rect 10919 5556 10931 5559
rect 11422 5556 11428 5568
rect 10919 5528 11428 5556
rect 10919 5525 10931 5528
rect 10873 5519 10931 5525
rect 11422 5516 11428 5528
rect 11480 5516 11486 5568
rect 1104 5466 13616 5488
rect 1104 5414 4078 5466
rect 4130 5414 4142 5466
rect 4194 5414 4206 5466
rect 4258 5414 4270 5466
rect 4322 5414 4334 5466
rect 4386 5414 7206 5466
rect 7258 5414 7270 5466
rect 7322 5414 7334 5466
rect 7386 5414 7398 5466
rect 7450 5414 7462 5466
rect 7514 5414 10334 5466
rect 10386 5414 10398 5466
rect 10450 5414 10462 5466
rect 10514 5414 10526 5466
rect 10578 5414 10590 5466
rect 10642 5414 13616 5466
rect 1104 5392 13616 5414
rect 3881 5355 3939 5361
rect 3881 5321 3893 5355
rect 3927 5352 3939 5355
rect 3970 5352 3976 5364
rect 3927 5324 3976 5352
rect 3927 5321 3939 5324
rect 3881 5315 3939 5321
rect 3970 5312 3976 5324
rect 4028 5312 4034 5364
rect 5534 5352 5540 5364
rect 4540 5324 5540 5352
rect 3878 5176 3884 5228
rect 3936 5216 3942 5228
rect 4540 5225 4568 5324
rect 5534 5312 5540 5324
rect 5592 5312 5598 5364
rect 8110 5352 8116 5364
rect 6886 5324 8116 5352
rect 4706 5244 4712 5296
rect 4764 5284 4770 5296
rect 4764 5256 5488 5284
rect 4764 5244 4770 5256
rect 4065 5219 4123 5225
rect 4065 5216 4077 5219
rect 3936 5188 4077 5216
rect 3936 5176 3942 5188
rect 4065 5185 4077 5188
rect 4111 5185 4123 5219
rect 4065 5179 4123 5185
rect 4341 5219 4399 5225
rect 4341 5185 4353 5219
rect 4387 5185 4399 5219
rect 4341 5179 4399 5185
rect 4525 5219 4583 5225
rect 4525 5185 4537 5219
rect 4571 5185 4583 5219
rect 5166 5216 5172 5228
rect 5127 5188 5172 5216
rect 4525 5179 4583 5185
rect 4356 5148 4384 5179
rect 5166 5176 5172 5188
rect 5224 5176 5230 5228
rect 5460 5225 5488 5256
rect 5445 5219 5503 5225
rect 5445 5185 5457 5219
rect 5491 5185 5503 5219
rect 5445 5179 5503 5185
rect 5629 5219 5687 5225
rect 5629 5185 5641 5219
rect 5675 5216 5687 5219
rect 6886 5216 6914 5324
rect 8110 5312 8116 5324
rect 8168 5352 8174 5364
rect 9582 5352 9588 5364
rect 8168 5324 9588 5352
rect 8168 5312 8174 5324
rect 9582 5312 9588 5324
rect 9640 5312 9646 5364
rect 10045 5355 10103 5361
rect 10045 5321 10057 5355
rect 10091 5352 10103 5355
rect 11330 5352 11336 5364
rect 10091 5324 11336 5352
rect 10091 5321 10103 5324
rect 10045 5315 10103 5321
rect 11330 5312 11336 5324
rect 11388 5312 11394 5364
rect 7469 5287 7527 5293
rect 7469 5253 7481 5287
rect 7515 5284 7527 5287
rect 7558 5284 7564 5296
rect 7515 5256 7564 5284
rect 7515 5253 7527 5256
rect 7469 5247 7527 5253
rect 7558 5244 7564 5256
rect 7616 5244 7622 5296
rect 9306 5244 9312 5296
rect 9364 5284 9370 5296
rect 9674 5284 9680 5296
rect 9364 5256 9680 5284
rect 9364 5244 9370 5256
rect 9674 5244 9680 5256
rect 9732 5284 9738 5296
rect 9732 5256 9904 5284
rect 9732 5244 9738 5256
rect 9401 5219 9459 5225
rect 5675 5188 6914 5216
rect 8602 5188 8800 5216
rect 5675 5185 5687 5188
rect 5629 5179 5687 5185
rect 4985 5151 5043 5157
rect 4985 5148 4997 5151
rect 4356 5120 4997 5148
rect 4985 5117 4997 5120
rect 5031 5117 5043 5151
rect 4985 5111 5043 5117
rect 7193 5151 7251 5157
rect 7193 5117 7205 5151
rect 7239 5148 7251 5151
rect 8662 5148 8668 5160
rect 7239 5120 8668 5148
rect 7239 5117 7251 5120
rect 7193 5111 7251 5117
rect 8662 5108 8668 5120
rect 8720 5108 8726 5160
rect 8772 5080 8800 5188
rect 9401 5185 9413 5219
rect 9447 5185 9459 5219
rect 9582 5216 9588 5228
rect 9543 5188 9588 5216
rect 9401 5179 9459 5185
rect 8941 5151 8999 5157
rect 8941 5117 8953 5151
rect 8987 5148 8999 5151
rect 9214 5148 9220 5160
rect 8987 5120 9220 5148
rect 8987 5117 8999 5120
rect 8941 5111 8999 5117
rect 9214 5108 9220 5120
rect 9272 5148 9278 5160
rect 9416 5148 9444 5179
rect 9582 5176 9588 5188
rect 9640 5176 9646 5228
rect 9876 5225 9904 5256
rect 9861 5219 9919 5225
rect 9861 5185 9873 5219
rect 9907 5185 9919 5219
rect 10686 5216 10692 5228
rect 10599 5188 10692 5216
rect 9861 5179 9919 5185
rect 10686 5176 10692 5188
rect 10744 5216 10750 5228
rect 12618 5216 12624 5228
rect 10744 5188 12624 5216
rect 10744 5176 10750 5188
rect 12618 5176 12624 5188
rect 12676 5176 12682 5228
rect 9272 5120 9444 5148
rect 9272 5108 9278 5120
rect 12710 5108 12716 5160
rect 12768 5148 12774 5160
rect 12897 5151 12955 5157
rect 12897 5148 12909 5151
rect 12768 5120 12909 5148
rect 12768 5108 12774 5120
rect 12897 5117 12909 5120
rect 12943 5117 12955 5151
rect 12897 5111 12955 5117
rect 8772 5052 10640 5080
rect 10612 5021 10640 5052
rect 10597 5015 10655 5021
rect 10597 4981 10609 5015
rect 10643 5012 10655 5015
rect 10778 5012 10784 5024
rect 10643 4984 10784 5012
rect 10643 4981 10655 4984
rect 10597 4975 10655 4981
rect 10778 4972 10784 4984
rect 10836 4972 10842 5024
rect 1104 4922 13616 4944
rect 1104 4870 2514 4922
rect 2566 4870 2578 4922
rect 2630 4870 2642 4922
rect 2694 4870 2706 4922
rect 2758 4870 2770 4922
rect 2822 4870 5642 4922
rect 5694 4870 5706 4922
rect 5758 4870 5770 4922
rect 5822 4870 5834 4922
rect 5886 4870 5898 4922
rect 5950 4870 8770 4922
rect 8822 4870 8834 4922
rect 8886 4870 8898 4922
rect 8950 4870 8962 4922
rect 9014 4870 9026 4922
rect 9078 4870 11898 4922
rect 11950 4870 11962 4922
rect 12014 4870 12026 4922
rect 12078 4870 12090 4922
rect 12142 4870 12154 4922
rect 12206 4870 13616 4922
rect 1104 4848 13616 4870
rect 6457 4675 6515 4681
rect 6457 4672 6469 4675
rect 3804 4644 6469 4672
rect 2130 4604 2136 4616
rect 2091 4576 2136 4604
rect 2130 4564 2136 4576
rect 2188 4564 2194 4616
rect 3234 4564 3240 4616
rect 3292 4604 3298 4616
rect 3804 4613 3832 4644
rect 6457 4641 6469 4644
rect 6503 4641 6515 4675
rect 6457 4635 6515 4641
rect 8662 4632 8668 4684
rect 8720 4672 8726 4684
rect 8941 4675 8999 4681
rect 8941 4672 8953 4675
rect 8720 4644 8953 4672
rect 8720 4632 8726 4644
rect 8941 4641 8953 4644
rect 8987 4641 8999 4675
rect 9214 4672 9220 4684
rect 9175 4644 9220 4672
rect 8941 4635 8999 4641
rect 9214 4632 9220 4644
rect 9272 4632 9278 4684
rect 11422 4672 11428 4684
rect 11383 4644 11428 4672
rect 11422 4632 11428 4644
rect 11480 4632 11486 4684
rect 3789 4607 3847 4613
rect 3789 4604 3801 4607
rect 3292 4576 3801 4604
rect 3292 4564 3298 4576
rect 3789 4573 3801 4576
rect 3835 4573 3847 4607
rect 3789 4567 3847 4573
rect 10226 4564 10232 4616
rect 10284 4604 10290 4616
rect 10686 4604 10692 4616
rect 10284 4576 10692 4604
rect 10284 4564 10290 4576
rect 10686 4564 10692 4576
rect 10744 4564 10750 4616
rect 11146 4604 11152 4616
rect 11107 4576 11152 4604
rect 11146 4564 11152 4576
rect 11204 4564 11210 4616
rect 5442 4496 5448 4548
rect 5500 4496 5506 4548
rect 6181 4539 6239 4545
rect 6181 4505 6193 4539
rect 6227 4536 6239 4539
rect 9214 4536 9220 4548
rect 6227 4508 9220 4536
rect 6227 4505 6239 4508
rect 6181 4499 6239 4505
rect 9214 4496 9220 4508
rect 9272 4496 9278 4548
rect 12710 4536 12716 4548
rect 12650 4508 12716 4536
rect 12710 4496 12716 4508
rect 12768 4496 12774 4548
rect 2317 4471 2375 4477
rect 2317 4437 2329 4471
rect 2363 4468 2375 4471
rect 2866 4468 2872 4480
rect 2363 4440 2872 4468
rect 2363 4437 2375 4440
rect 2317 4431 2375 4437
rect 2866 4428 2872 4440
rect 2924 4428 2930 4480
rect 3786 4428 3792 4480
rect 3844 4468 3850 4480
rect 3973 4471 4031 4477
rect 3973 4468 3985 4471
rect 3844 4440 3985 4468
rect 3844 4428 3850 4440
rect 3973 4437 3985 4440
rect 4019 4437 4031 4471
rect 4706 4468 4712 4480
rect 4667 4440 4712 4468
rect 3973 4431 4031 4437
rect 4706 4428 4712 4440
rect 4764 4428 4770 4480
rect 10686 4468 10692 4480
rect 10647 4440 10692 4468
rect 10686 4428 10692 4440
rect 10744 4428 10750 4480
rect 12802 4428 12808 4480
rect 12860 4468 12866 4480
rect 12897 4471 12955 4477
rect 12897 4468 12909 4471
rect 12860 4440 12909 4468
rect 12860 4428 12866 4440
rect 12897 4437 12909 4440
rect 12943 4437 12955 4471
rect 12897 4431 12955 4437
rect 1104 4378 13616 4400
rect 1104 4326 4078 4378
rect 4130 4326 4142 4378
rect 4194 4326 4206 4378
rect 4258 4326 4270 4378
rect 4322 4326 4334 4378
rect 4386 4326 7206 4378
rect 7258 4326 7270 4378
rect 7322 4326 7334 4378
rect 7386 4326 7398 4378
rect 7450 4326 7462 4378
rect 7514 4326 10334 4378
rect 10386 4326 10398 4378
rect 10450 4326 10462 4378
rect 10514 4326 10526 4378
rect 10578 4326 10590 4378
rect 10642 4326 13616 4378
rect 1104 4304 13616 4326
rect 2130 4224 2136 4276
rect 2188 4264 2194 4276
rect 2685 4267 2743 4273
rect 2685 4264 2697 4267
rect 2188 4236 2697 4264
rect 2188 4224 2194 4236
rect 2685 4233 2697 4236
rect 2731 4233 2743 4267
rect 2685 4227 2743 4233
rect 4985 4267 5043 4273
rect 4985 4233 4997 4267
rect 5031 4264 5043 4267
rect 5166 4264 5172 4276
rect 5031 4236 5172 4264
rect 5031 4233 5043 4236
rect 4985 4227 5043 4233
rect 5166 4224 5172 4236
rect 5224 4224 5230 4276
rect 9214 4264 9220 4276
rect 9175 4236 9220 4264
rect 9214 4224 9220 4236
rect 9272 4224 9278 4276
rect 11146 4264 11152 4276
rect 9416 4236 11152 4264
rect 5442 4196 5448 4208
rect 4738 4168 5448 4196
rect 5442 4156 5448 4168
rect 5500 4156 5506 4208
rect 6917 4199 6975 4205
rect 6917 4165 6929 4199
rect 6963 4196 6975 4199
rect 7558 4196 7564 4208
rect 6963 4168 7564 4196
rect 6963 4165 6975 4168
rect 6917 4159 6975 4165
rect 7558 4156 7564 4168
rect 7616 4156 7622 4208
rect 8662 4156 8668 4208
rect 8720 4196 8726 4208
rect 9416 4196 9444 4236
rect 8720 4168 9444 4196
rect 8720 4156 8726 4168
rect 10226 4156 10232 4208
rect 10284 4156 10290 4208
rect 10686 4196 10692 4208
rect 10647 4168 10692 4196
rect 10686 4156 10692 4168
rect 10744 4156 10750 4208
rect 10888 4196 10916 4236
rect 11146 4224 11152 4236
rect 11204 4224 11210 4276
rect 12710 4264 12716 4276
rect 12671 4236 12716 4264
rect 12710 4224 12716 4236
rect 12768 4224 12774 4276
rect 10888 4168 11008 4196
rect 2314 4128 2320 4140
rect 2275 4100 2320 4128
rect 2314 4088 2320 4100
rect 2372 4088 2378 4140
rect 3234 4128 3240 4140
rect 3195 4100 3240 4128
rect 3234 4088 3240 4100
rect 3292 4088 3298 4140
rect 7006 4088 7012 4140
rect 7064 4128 7070 4140
rect 8110 4128 8116 4140
rect 7064 4100 7109 4128
rect 8071 4100 8116 4128
rect 7064 4088 7070 4100
rect 8110 4088 8116 4100
rect 8168 4088 8174 4140
rect 8297 4131 8355 4137
rect 8297 4097 8309 4131
rect 8343 4097 8355 4131
rect 8570 4128 8576 4140
rect 8531 4100 8576 4128
rect 8297 4091 8355 4097
rect 2133 4063 2191 4069
rect 2133 4029 2145 4063
rect 2179 4029 2191 4063
rect 2133 4023 2191 4029
rect 2225 4063 2283 4069
rect 2225 4029 2237 4063
rect 2271 4060 2283 4063
rect 3142 4060 3148 4072
rect 2271 4032 3148 4060
rect 2271 4029 2283 4032
rect 2225 4023 2283 4029
rect 2148 3924 2176 4023
rect 3142 4020 3148 4032
rect 3200 4020 3206 4072
rect 3510 4060 3516 4072
rect 3471 4032 3516 4060
rect 3510 4020 3516 4032
rect 3568 4020 3574 4072
rect 7101 4063 7159 4069
rect 7101 4060 7113 4063
rect 6886 4032 7113 4060
rect 6886 3992 6914 4032
rect 7101 4029 7113 4032
rect 7147 4029 7159 4063
rect 8312 4060 8340 4091
rect 8570 4088 8576 4100
rect 8628 4088 8634 4140
rect 10980 4137 11008 4168
rect 10965 4131 11023 4137
rect 10965 4097 10977 4131
rect 11011 4097 11023 4131
rect 12894 4128 12900 4140
rect 12855 4100 12900 4128
rect 10965 4091 11023 4097
rect 12894 4088 12900 4100
rect 12952 4088 12958 4140
rect 10686 4060 10692 4072
rect 8312 4032 10692 4060
rect 7101 4023 7159 4029
rect 10686 4020 10692 4032
rect 10744 4020 10750 4072
rect 4540 3964 6914 3992
rect 2406 3924 2412 3936
rect 2148 3896 2412 3924
rect 2406 3884 2412 3896
rect 2464 3924 2470 3936
rect 4540 3924 4568 3964
rect 6546 3924 6552 3936
rect 2464 3896 4568 3924
rect 6507 3896 6552 3924
rect 2464 3884 2470 3896
rect 6546 3884 6552 3896
rect 6604 3884 6610 3936
rect 8662 3884 8668 3936
rect 8720 3924 8726 3936
rect 8757 3927 8815 3933
rect 8757 3924 8769 3927
rect 8720 3896 8769 3924
rect 8720 3884 8726 3896
rect 8757 3893 8769 3896
rect 8803 3893 8815 3927
rect 8757 3887 8815 3893
rect 1104 3834 13616 3856
rect 1104 3782 2514 3834
rect 2566 3782 2578 3834
rect 2630 3782 2642 3834
rect 2694 3782 2706 3834
rect 2758 3782 2770 3834
rect 2822 3782 5642 3834
rect 5694 3782 5706 3834
rect 5758 3782 5770 3834
rect 5822 3782 5834 3834
rect 5886 3782 5898 3834
rect 5950 3782 8770 3834
rect 8822 3782 8834 3834
rect 8886 3782 8898 3834
rect 8950 3782 8962 3834
rect 9014 3782 9026 3834
rect 9078 3782 11898 3834
rect 11950 3782 11962 3834
rect 12014 3782 12026 3834
rect 12078 3782 12090 3834
rect 12142 3782 12154 3834
rect 12206 3782 13616 3834
rect 1104 3760 13616 3782
rect 1397 3723 1455 3729
rect 1397 3689 1409 3723
rect 1443 3720 1455 3723
rect 1670 3720 1676 3732
rect 1443 3692 1676 3720
rect 1443 3689 1455 3692
rect 1397 3683 1455 3689
rect 1670 3680 1676 3692
rect 1728 3720 1734 3732
rect 2314 3720 2320 3732
rect 1728 3692 2320 3720
rect 1728 3680 1734 3692
rect 2314 3680 2320 3692
rect 2372 3680 2378 3732
rect 3602 3680 3608 3732
rect 3660 3720 3666 3732
rect 3973 3723 4031 3729
rect 3973 3720 3985 3723
rect 3660 3692 3985 3720
rect 3660 3680 3666 3692
rect 3973 3689 3985 3692
rect 4019 3689 4031 3723
rect 7558 3720 7564 3732
rect 7519 3692 7564 3720
rect 3973 3683 4031 3689
rect 7558 3680 7564 3692
rect 7616 3680 7622 3732
rect 8389 3723 8447 3729
rect 8389 3689 8401 3723
rect 8435 3720 8447 3723
rect 8570 3720 8576 3732
rect 8435 3692 8576 3720
rect 8435 3689 8447 3692
rect 8389 3683 8447 3689
rect 8570 3680 8576 3692
rect 8628 3680 8634 3732
rect 10686 3720 10692 3732
rect 10647 3692 10692 3720
rect 10686 3680 10692 3692
rect 10744 3680 10750 3732
rect 2866 3584 2872 3596
rect 2827 3556 2872 3584
rect 2866 3544 2872 3556
rect 2924 3544 2930 3596
rect 5828 3556 8248 3584
rect 3145 3519 3203 3525
rect 3145 3485 3157 3519
rect 3191 3516 3203 3519
rect 3786 3516 3792 3528
rect 3191 3488 3792 3516
rect 3191 3485 3203 3488
rect 3145 3479 3203 3485
rect 3786 3476 3792 3488
rect 3844 3476 3850 3528
rect 5442 3476 5448 3528
rect 5500 3516 5506 3528
rect 5828 3525 5856 3556
rect 8220 3525 8248 3556
rect 8662 3544 8668 3596
rect 8720 3584 8726 3596
rect 9217 3587 9275 3593
rect 9217 3584 9229 3587
rect 8720 3556 9229 3584
rect 8720 3544 8726 3556
rect 9217 3553 9229 3556
rect 9263 3553 9275 3587
rect 9217 3547 9275 3553
rect 5813 3519 5871 3525
rect 5813 3516 5825 3519
rect 5500 3488 5825 3516
rect 5500 3476 5506 3488
rect 5813 3485 5825 3488
rect 5859 3485 5871 3519
rect 5813 3479 5871 3485
rect 8205 3519 8263 3525
rect 8205 3485 8217 3519
rect 8251 3516 8263 3519
rect 8941 3519 8999 3525
rect 8941 3516 8953 3519
rect 8251 3488 8953 3516
rect 8251 3485 8263 3488
rect 8205 3479 8263 3485
rect 8941 3485 8953 3488
rect 8987 3485 8999 3519
rect 8941 3479 8999 3485
rect 3418 3448 3424 3460
rect 2438 3420 3424 3448
rect 3418 3408 3424 3420
rect 3476 3408 3482 3460
rect 6089 3451 6147 3457
rect 6089 3417 6101 3451
rect 6135 3448 6147 3451
rect 6362 3448 6368 3460
rect 6135 3420 6368 3448
rect 6135 3417 6147 3420
rect 6089 3411 6147 3417
rect 6362 3408 6368 3420
rect 6420 3408 6426 3460
rect 10778 3448 10784 3460
rect 7314 3420 8156 3448
rect 10442 3420 10784 3448
rect 7098 3340 7104 3392
rect 7156 3380 7162 3392
rect 7392 3380 7420 3420
rect 7156 3352 7420 3380
rect 8128 3380 8156 3420
rect 10520 3380 10548 3420
rect 10778 3408 10784 3420
rect 10836 3408 10842 3460
rect 8128 3352 10548 3380
rect 7156 3340 7162 3352
rect 1104 3290 13616 3312
rect 1104 3238 4078 3290
rect 4130 3238 4142 3290
rect 4194 3238 4206 3290
rect 4258 3238 4270 3290
rect 4322 3238 4334 3290
rect 4386 3238 7206 3290
rect 7258 3238 7270 3290
rect 7322 3238 7334 3290
rect 7386 3238 7398 3290
rect 7450 3238 7462 3290
rect 7514 3238 10334 3290
rect 10386 3238 10398 3290
rect 10450 3238 10462 3290
rect 10514 3238 10526 3290
rect 10578 3238 10590 3290
rect 10642 3238 13616 3290
rect 1104 3216 13616 3238
rect 1486 3176 1492 3188
rect 1447 3148 1492 3176
rect 1486 3136 1492 3148
rect 1544 3136 1550 3188
rect 2409 3179 2467 3185
rect 2409 3145 2421 3179
rect 2455 3176 2467 3179
rect 3510 3176 3516 3188
rect 2455 3148 3516 3176
rect 2455 3145 2467 3148
rect 2409 3139 2467 3145
rect 3510 3136 3516 3148
rect 3568 3136 3574 3188
rect 6362 3176 6368 3188
rect 3712 3148 5396 3176
rect 6323 3148 6368 3176
rect 3418 3068 3424 3120
rect 3476 3108 3482 3120
rect 3712 3108 3740 3148
rect 5368 3120 5396 3148
rect 6362 3136 6368 3148
rect 6420 3136 6426 3188
rect 3476 3080 3740 3108
rect 3476 3068 3482 3080
rect 3786 3068 3792 3120
rect 3844 3108 3850 3120
rect 3844 3080 4200 3108
rect 3844 3068 3850 3080
rect 1670 3040 1676 3052
rect 1631 3012 1676 3040
rect 1670 3000 1676 3012
rect 1728 3000 1734 3052
rect 4172 3049 4200 3080
rect 5350 3068 5356 3120
rect 5408 3108 5414 3120
rect 7009 3111 7067 3117
rect 7009 3108 7021 3111
rect 5408 3080 7021 3108
rect 5408 3068 5414 3080
rect 7009 3077 7021 3080
rect 7055 3077 7067 3111
rect 7009 3071 7067 3077
rect 7098 3068 7104 3120
rect 7156 3108 7162 3120
rect 7193 3111 7251 3117
rect 7193 3108 7205 3111
rect 7156 3080 7205 3108
rect 7156 3068 7162 3080
rect 7193 3077 7205 3080
rect 7239 3077 7251 3111
rect 7193 3071 7251 3077
rect 4157 3043 4215 3049
rect 4157 3009 4169 3043
rect 4203 3009 4215 3043
rect 6546 3040 6552 3052
rect 6507 3012 6552 3040
rect 4157 3003 4215 3009
rect 6546 3000 6552 3012
rect 6604 3000 6610 3052
rect 3881 2975 3939 2981
rect 3881 2941 3893 2975
rect 3927 2972 3939 2975
rect 4706 2972 4712 2984
rect 3927 2944 4712 2972
rect 3927 2941 3939 2944
rect 3881 2935 3939 2941
rect 4706 2932 4712 2944
rect 4764 2932 4770 2984
rect 1104 2746 13616 2768
rect 1104 2694 2514 2746
rect 2566 2694 2578 2746
rect 2630 2694 2642 2746
rect 2694 2694 2706 2746
rect 2758 2694 2770 2746
rect 2822 2694 5642 2746
rect 5694 2694 5706 2746
rect 5758 2694 5770 2746
rect 5822 2694 5834 2746
rect 5886 2694 5898 2746
rect 5950 2694 8770 2746
rect 8822 2694 8834 2746
rect 8886 2694 8898 2746
rect 8950 2694 8962 2746
rect 9014 2694 9026 2746
rect 9078 2694 11898 2746
rect 11950 2694 11962 2746
rect 12014 2694 12026 2746
rect 12078 2694 12090 2746
rect 12142 2694 12154 2746
rect 12206 2694 13616 2746
rect 1104 2672 13616 2694
rect 3237 2635 3295 2641
rect 3237 2601 3249 2635
rect 3283 2632 3295 2635
rect 5442 2632 5448 2644
rect 3283 2604 5448 2632
rect 3283 2601 3295 2604
rect 3237 2595 3295 2601
rect 5442 2592 5448 2604
rect 5500 2592 5506 2644
rect 2041 2567 2099 2573
rect 2041 2533 2053 2567
rect 2087 2564 2099 2567
rect 4430 2564 4436 2576
rect 2087 2536 4436 2564
rect 2087 2533 2099 2536
rect 2041 2527 2099 2533
rect 4430 2524 4436 2536
rect 4488 2524 4494 2576
rect 3234 2456 3240 2508
rect 3292 2496 3298 2508
rect 4341 2499 4399 2505
rect 4341 2496 4353 2499
rect 3292 2468 4353 2496
rect 3292 2456 3298 2468
rect 4341 2465 4353 2468
rect 4387 2465 4399 2499
rect 4341 2459 4399 2465
rect 3053 2431 3111 2437
rect 3053 2397 3065 2431
rect 3099 2428 3111 2431
rect 3252 2428 3280 2456
rect 3099 2400 3280 2428
rect 3099 2397 3111 2400
rect 3053 2391 3111 2397
rect 3878 2388 3884 2440
rect 3936 2428 3942 2440
rect 4065 2431 4123 2437
rect 4065 2428 4077 2431
rect 3936 2400 4077 2428
rect 3936 2388 3942 2400
rect 4065 2397 4077 2400
rect 4111 2397 4123 2431
rect 4065 2391 4123 2397
rect 7558 2388 7564 2440
rect 7616 2428 7622 2440
rect 7837 2431 7895 2437
rect 7837 2428 7849 2431
rect 7616 2400 7849 2428
rect 7616 2388 7622 2400
rect 7837 2397 7849 2400
rect 7883 2397 7895 2431
rect 7837 2391 7895 2397
rect 10686 2388 10692 2440
rect 10744 2428 10750 2440
rect 11701 2431 11759 2437
rect 11701 2428 11713 2431
rect 10744 2400 11713 2428
rect 10744 2388 10750 2400
rect 11701 2397 11713 2400
rect 11747 2397 11759 2431
rect 11701 2391 11759 2397
rect 12621 2431 12679 2437
rect 12621 2397 12633 2431
rect 12667 2428 12679 2431
rect 12802 2428 12808 2440
rect 12667 2400 12808 2428
rect 12667 2397 12679 2400
rect 12621 2391 12679 2397
rect 12802 2388 12808 2400
rect 12860 2388 12866 2440
rect 14 2320 20 2372
rect 72 2360 78 2372
rect 1857 2363 1915 2369
rect 1857 2360 1869 2363
rect 72 2332 1869 2360
rect 72 2320 78 2332
rect 1857 2329 1869 2332
rect 1903 2329 1915 2363
rect 1857 2323 1915 2329
rect 7742 2252 7748 2304
rect 7800 2292 7806 2304
rect 8021 2295 8079 2301
rect 8021 2292 8033 2295
rect 7800 2264 8033 2292
rect 7800 2252 7806 2264
rect 8021 2261 8033 2264
rect 8067 2261 8079 2295
rect 8021 2255 8079 2261
rect 11606 2252 11612 2304
rect 11664 2292 11670 2304
rect 11885 2295 11943 2301
rect 11885 2292 11897 2295
rect 11664 2264 11897 2292
rect 11664 2252 11670 2264
rect 11885 2261 11897 2264
rect 11931 2261 11943 2295
rect 11885 2255 11943 2261
rect 12342 2252 12348 2304
rect 12400 2292 12406 2304
rect 12805 2295 12863 2301
rect 12805 2292 12817 2295
rect 12400 2264 12817 2292
rect 12400 2252 12406 2264
rect 12805 2261 12817 2264
rect 12851 2261 12863 2295
rect 12805 2255 12863 2261
rect 1104 2202 13616 2224
rect 1104 2150 4078 2202
rect 4130 2150 4142 2202
rect 4194 2150 4206 2202
rect 4258 2150 4270 2202
rect 4322 2150 4334 2202
rect 4386 2150 7206 2202
rect 7258 2150 7270 2202
rect 7322 2150 7334 2202
rect 7386 2150 7398 2202
rect 7450 2150 7462 2202
rect 7514 2150 10334 2202
rect 10386 2150 10398 2202
rect 10450 2150 10462 2202
rect 10514 2150 10526 2202
rect 10578 2150 10590 2202
rect 10642 2150 13616 2202
rect 1104 2128 13616 2150
<< via1 >>
rect 2514 14662 2566 14714
rect 2578 14662 2630 14714
rect 2642 14662 2694 14714
rect 2706 14662 2758 14714
rect 2770 14662 2822 14714
rect 5642 14662 5694 14714
rect 5706 14662 5758 14714
rect 5770 14662 5822 14714
rect 5834 14662 5886 14714
rect 5898 14662 5950 14714
rect 8770 14662 8822 14714
rect 8834 14662 8886 14714
rect 8898 14662 8950 14714
rect 8962 14662 9014 14714
rect 9026 14662 9078 14714
rect 11898 14662 11950 14714
rect 11962 14662 12014 14714
rect 12026 14662 12078 14714
rect 12090 14662 12142 14714
rect 12154 14662 12206 14714
rect 1492 14603 1544 14612
rect 1492 14569 1501 14603
rect 1501 14569 1535 14603
rect 1535 14569 1544 14603
rect 1492 14560 1544 14569
rect 6460 14560 6512 14612
rect 10324 14560 10376 14612
rect 14188 14560 14240 14612
rect 2412 14356 2464 14408
rect 7012 14356 7064 14408
rect 10692 14399 10744 14408
rect 10692 14365 10701 14399
rect 10701 14365 10735 14399
rect 10735 14365 10744 14399
rect 10692 14356 10744 14365
rect 12440 14356 12492 14408
rect 3240 14288 3292 14340
rect 4988 14220 5040 14272
rect 4078 14118 4130 14170
rect 4142 14118 4194 14170
rect 4206 14118 4258 14170
rect 4270 14118 4322 14170
rect 4334 14118 4386 14170
rect 7206 14118 7258 14170
rect 7270 14118 7322 14170
rect 7334 14118 7386 14170
rect 7398 14118 7450 14170
rect 7462 14118 7514 14170
rect 10334 14118 10386 14170
rect 10398 14118 10450 14170
rect 10462 14118 10514 14170
rect 10526 14118 10578 14170
rect 10590 14118 10642 14170
rect 6368 13923 6420 13932
rect 6368 13889 6377 13923
rect 6377 13889 6411 13923
rect 6411 13889 6420 13923
rect 6368 13880 6420 13889
rect 9772 13880 9824 13932
rect 10232 13923 10284 13932
rect 10232 13889 10241 13923
rect 10241 13889 10275 13923
rect 10275 13889 10284 13923
rect 10232 13880 10284 13889
rect 10048 13855 10100 13864
rect 10048 13821 10057 13855
rect 10057 13821 10091 13855
rect 10091 13821 10100 13855
rect 10048 13812 10100 13821
rect 4252 13719 4304 13728
rect 4252 13685 4261 13719
rect 4261 13685 4295 13719
rect 4295 13685 4304 13719
rect 4252 13676 4304 13685
rect 6828 13676 6880 13728
rect 9220 13719 9272 13728
rect 9220 13685 9229 13719
rect 9229 13685 9263 13719
rect 9263 13685 9272 13719
rect 9220 13676 9272 13685
rect 2514 13574 2566 13626
rect 2578 13574 2630 13626
rect 2642 13574 2694 13626
rect 2706 13574 2758 13626
rect 2770 13574 2822 13626
rect 5642 13574 5694 13626
rect 5706 13574 5758 13626
rect 5770 13574 5822 13626
rect 5834 13574 5886 13626
rect 5898 13574 5950 13626
rect 8770 13574 8822 13626
rect 8834 13574 8886 13626
rect 8898 13574 8950 13626
rect 8962 13574 9014 13626
rect 9026 13574 9078 13626
rect 11898 13574 11950 13626
rect 11962 13574 12014 13626
rect 12026 13574 12078 13626
rect 12090 13574 12142 13626
rect 12154 13574 12206 13626
rect 10692 13515 10744 13524
rect 10692 13481 10701 13515
rect 10701 13481 10735 13515
rect 10735 13481 10744 13515
rect 10692 13472 10744 13481
rect 4252 13379 4304 13388
rect 4252 13345 4261 13379
rect 4261 13345 4295 13379
rect 4295 13345 4304 13379
rect 4252 13336 4304 13345
rect 6828 13379 6880 13388
rect 6828 13345 6837 13379
rect 6837 13345 6871 13379
rect 6871 13345 6880 13379
rect 6828 13336 6880 13345
rect 9220 13379 9272 13388
rect 9220 13345 9229 13379
rect 9229 13345 9263 13379
rect 9263 13345 9272 13379
rect 9220 13336 9272 13345
rect 4344 13268 4396 13320
rect 6552 13311 6604 13320
rect 6552 13277 6561 13311
rect 6561 13277 6595 13311
rect 6595 13277 6604 13311
rect 6552 13268 6604 13277
rect 5448 13132 5500 13184
rect 8208 13200 8260 13252
rect 12992 13268 13044 13320
rect 10968 13200 11020 13252
rect 8300 13175 8352 13184
rect 8300 13141 8309 13175
rect 8309 13141 8343 13175
rect 8343 13141 8352 13175
rect 8300 13132 8352 13141
rect 9588 13132 9640 13184
rect 12808 13175 12860 13184
rect 12808 13141 12817 13175
rect 12817 13141 12851 13175
rect 12851 13141 12860 13175
rect 12808 13132 12860 13141
rect 4078 13030 4130 13082
rect 4142 13030 4194 13082
rect 4206 13030 4258 13082
rect 4270 13030 4322 13082
rect 4334 13030 4386 13082
rect 7206 13030 7258 13082
rect 7270 13030 7322 13082
rect 7334 13030 7386 13082
rect 7398 13030 7450 13082
rect 7462 13030 7514 13082
rect 10334 13030 10386 13082
rect 10398 13030 10450 13082
rect 10462 13030 10514 13082
rect 10526 13030 10578 13082
rect 10590 13030 10642 13082
rect 6368 12928 6420 12980
rect 9772 12928 9824 12980
rect 10692 12928 10744 12980
rect 4988 12835 5040 12844
rect 4988 12801 4997 12835
rect 4997 12801 5031 12835
rect 5031 12801 5040 12835
rect 4988 12792 5040 12801
rect 5264 12835 5316 12844
rect 5264 12801 5273 12835
rect 5273 12801 5307 12835
rect 5307 12801 5316 12835
rect 5264 12792 5316 12801
rect 5448 12792 5500 12844
rect 12716 12792 12768 12844
rect 10140 12767 10192 12776
rect 10140 12733 10149 12767
rect 10149 12733 10183 12767
rect 10183 12733 10192 12767
rect 10140 12724 10192 12733
rect 10232 12767 10284 12776
rect 10232 12733 10241 12767
rect 10241 12733 10275 12767
rect 10275 12733 10284 12767
rect 10232 12724 10284 12733
rect 12808 12724 12860 12776
rect 6276 12656 6328 12708
rect 10968 12656 11020 12708
rect 4896 12588 4948 12640
rect 2514 12486 2566 12538
rect 2578 12486 2630 12538
rect 2642 12486 2694 12538
rect 2706 12486 2758 12538
rect 2770 12486 2822 12538
rect 5642 12486 5694 12538
rect 5706 12486 5758 12538
rect 5770 12486 5822 12538
rect 5834 12486 5886 12538
rect 5898 12486 5950 12538
rect 8770 12486 8822 12538
rect 8834 12486 8886 12538
rect 8898 12486 8950 12538
rect 8962 12486 9014 12538
rect 9026 12486 9078 12538
rect 11898 12486 11950 12538
rect 11962 12486 12014 12538
rect 12026 12486 12078 12538
rect 12090 12486 12142 12538
rect 12154 12486 12206 12538
rect 6276 12384 6328 12436
rect 4436 12248 4488 12300
rect 4620 12291 4672 12300
rect 4620 12257 4629 12291
rect 4629 12257 4663 12291
rect 4663 12257 4672 12291
rect 4620 12248 4672 12257
rect 4896 12291 4948 12300
rect 4896 12257 4905 12291
rect 4905 12257 4939 12291
rect 4939 12257 4948 12291
rect 4896 12248 4948 12257
rect 9588 12223 9640 12232
rect 9588 12189 9597 12223
rect 9597 12189 9631 12223
rect 9631 12189 9640 12223
rect 9588 12180 9640 12189
rect 10968 12180 11020 12232
rect 8208 12112 8260 12164
rect 9128 12112 9180 12164
rect 7932 12044 7984 12096
rect 10048 12044 10100 12096
rect 11336 12087 11388 12096
rect 11336 12053 11345 12087
rect 11345 12053 11379 12087
rect 11379 12053 11388 12087
rect 11336 12044 11388 12053
rect 4078 11942 4130 11994
rect 4142 11942 4194 11994
rect 4206 11942 4258 11994
rect 4270 11942 4322 11994
rect 4334 11942 4386 11994
rect 7206 11942 7258 11994
rect 7270 11942 7322 11994
rect 7334 11942 7386 11994
rect 7398 11942 7450 11994
rect 7462 11942 7514 11994
rect 10334 11942 10386 11994
rect 10398 11942 10450 11994
rect 10462 11942 10514 11994
rect 10526 11942 10578 11994
rect 10590 11942 10642 11994
rect 9128 11840 9180 11892
rect 2412 11772 2464 11824
rect 2964 11772 3016 11824
rect 9680 11772 9732 11824
rect 10968 11772 11020 11824
rect 2044 11704 2096 11756
rect 6552 11704 6604 11756
rect 2320 11636 2372 11688
rect 4160 11679 4212 11688
rect 4160 11645 4169 11679
rect 4169 11645 4203 11679
rect 4203 11645 4212 11679
rect 4160 11636 4212 11645
rect 5264 11636 5316 11688
rect 1492 11611 1544 11620
rect 1492 11577 1501 11611
rect 1501 11577 1535 11611
rect 1535 11577 1544 11611
rect 1492 11568 1544 11577
rect 8392 11636 8444 11688
rect 2412 11500 2464 11552
rect 7932 11500 7984 11552
rect 9588 11500 9640 11552
rect 2514 11398 2566 11450
rect 2578 11398 2630 11450
rect 2642 11398 2694 11450
rect 2706 11398 2758 11450
rect 2770 11398 2822 11450
rect 5642 11398 5694 11450
rect 5706 11398 5758 11450
rect 5770 11398 5822 11450
rect 5834 11398 5886 11450
rect 5898 11398 5950 11450
rect 8770 11398 8822 11450
rect 8834 11398 8886 11450
rect 8898 11398 8950 11450
rect 8962 11398 9014 11450
rect 9026 11398 9078 11450
rect 11898 11398 11950 11450
rect 11962 11398 12014 11450
rect 12026 11398 12078 11450
rect 12090 11398 12142 11450
rect 12154 11398 12206 11450
rect 8392 11339 8444 11348
rect 8392 11305 8401 11339
rect 8401 11305 8435 11339
rect 8435 11305 8444 11339
rect 8392 11296 8444 11305
rect 12808 11339 12860 11348
rect 12808 11305 12817 11339
rect 12817 11305 12851 11339
rect 12851 11305 12860 11339
rect 12808 11296 12860 11305
rect 6552 11160 6604 11212
rect 9588 11160 9640 11212
rect 11336 11203 11388 11212
rect 11336 11169 11345 11203
rect 11345 11169 11379 11203
rect 11379 11169 11388 11203
rect 11336 11160 11388 11169
rect 4160 11092 4212 11144
rect 4436 11135 4488 11144
rect 2044 11024 2096 11076
rect 4436 11101 4445 11135
rect 4445 11101 4479 11135
rect 4479 11101 4488 11135
rect 4436 11092 4488 11101
rect 9680 11092 9732 11144
rect 6920 11067 6972 11076
rect 6920 11033 6929 11067
rect 6929 11033 6963 11067
rect 6963 11033 6972 11067
rect 6920 11024 6972 11033
rect 8208 11024 8260 11076
rect 12716 11024 12768 11076
rect 3792 10999 3844 11008
rect 3792 10965 3801 10999
rect 3801 10965 3835 10999
rect 3835 10965 3844 10999
rect 3792 10956 3844 10965
rect 4078 10854 4130 10906
rect 4142 10854 4194 10906
rect 4206 10854 4258 10906
rect 4270 10854 4322 10906
rect 4334 10854 4386 10906
rect 7206 10854 7258 10906
rect 7270 10854 7322 10906
rect 7334 10854 7386 10906
rect 7398 10854 7450 10906
rect 7462 10854 7514 10906
rect 10334 10854 10386 10906
rect 10398 10854 10450 10906
rect 10462 10854 10514 10906
rect 10526 10854 10578 10906
rect 10590 10854 10642 10906
rect 2044 10795 2096 10804
rect 2044 10761 2053 10795
rect 2053 10761 2087 10795
rect 2087 10761 2096 10795
rect 2044 10752 2096 10761
rect 2872 10684 2924 10736
rect 3792 10684 3844 10736
rect 8300 10684 8352 10736
rect 10140 10684 10192 10736
rect 9128 10659 9180 10668
rect 1400 10548 1452 10600
rect 2320 10548 2372 10600
rect 7656 10548 7708 10600
rect 9128 10625 9137 10659
rect 9137 10625 9171 10659
rect 9171 10625 9180 10659
rect 9128 10616 9180 10625
rect 9956 10659 10008 10668
rect 9956 10625 9965 10659
rect 9965 10625 9999 10659
rect 9999 10625 10008 10659
rect 9956 10616 10008 10625
rect 10416 10659 10468 10668
rect 10416 10625 10425 10659
rect 10425 10625 10459 10659
rect 10459 10625 10468 10659
rect 10416 10616 10468 10625
rect 8116 10412 8168 10464
rect 9772 10455 9824 10464
rect 9772 10421 9781 10455
rect 9781 10421 9815 10455
rect 9815 10421 9824 10455
rect 9772 10412 9824 10421
rect 2514 10310 2566 10362
rect 2578 10310 2630 10362
rect 2642 10310 2694 10362
rect 2706 10310 2758 10362
rect 2770 10310 2822 10362
rect 5642 10310 5694 10362
rect 5706 10310 5758 10362
rect 5770 10310 5822 10362
rect 5834 10310 5886 10362
rect 5898 10310 5950 10362
rect 8770 10310 8822 10362
rect 8834 10310 8886 10362
rect 8898 10310 8950 10362
rect 8962 10310 9014 10362
rect 9026 10310 9078 10362
rect 11898 10310 11950 10362
rect 11962 10310 12014 10362
rect 12026 10310 12078 10362
rect 12090 10310 12142 10362
rect 12154 10310 12206 10362
rect 6276 10208 6328 10260
rect 6920 10208 6972 10260
rect 7656 10251 7708 10260
rect 7656 10217 7665 10251
rect 7665 10217 7699 10251
rect 7699 10217 7708 10251
rect 7656 10208 7708 10217
rect 4436 10072 4488 10124
rect 8116 10072 8168 10124
rect 9772 10115 9824 10124
rect 9772 10081 9781 10115
rect 9781 10081 9815 10115
rect 9815 10081 9824 10115
rect 9772 10072 9824 10081
rect 10416 10072 10468 10124
rect 12624 10072 12676 10124
rect 12808 10072 12860 10124
rect 4620 10004 4672 10056
rect 4988 10047 5040 10056
rect 4988 10013 4997 10047
rect 4997 10013 5031 10047
rect 5031 10013 5040 10047
rect 4988 10004 5040 10013
rect 9496 10047 9548 10056
rect 9496 10013 9505 10047
rect 9505 10013 9539 10047
rect 9539 10013 9548 10047
rect 9496 10004 9548 10013
rect 12440 10047 12492 10056
rect 12440 10013 12449 10047
rect 12449 10013 12483 10047
rect 12483 10013 12492 10047
rect 12440 10004 12492 10013
rect 3056 9868 3108 9920
rect 4528 9868 4580 9920
rect 6276 9936 6328 9988
rect 6920 9936 6972 9988
rect 12716 9936 12768 9988
rect 6552 9868 6604 9920
rect 12164 9868 12216 9920
rect 12532 9911 12584 9920
rect 12532 9877 12541 9911
rect 12541 9877 12575 9911
rect 12575 9877 12584 9911
rect 12532 9868 12584 9877
rect 4078 9766 4130 9818
rect 4142 9766 4194 9818
rect 4206 9766 4258 9818
rect 4270 9766 4322 9818
rect 4334 9766 4386 9818
rect 7206 9766 7258 9818
rect 7270 9766 7322 9818
rect 7334 9766 7386 9818
rect 7398 9766 7450 9818
rect 7462 9766 7514 9818
rect 10334 9766 10386 9818
rect 10398 9766 10450 9818
rect 10462 9766 10514 9818
rect 10526 9766 10578 9818
rect 10590 9766 10642 9818
rect 4528 9596 4580 9648
rect 2872 9528 2924 9580
rect 1400 9460 1452 9512
rect 1768 9503 1820 9512
rect 1768 9469 1777 9503
rect 1777 9469 1811 9503
rect 1811 9469 1820 9503
rect 1768 9460 1820 9469
rect 3240 9503 3292 9512
rect 3240 9469 3249 9503
rect 3249 9469 3283 9503
rect 3283 9469 3292 9503
rect 3240 9460 3292 9469
rect 3976 9503 4028 9512
rect 3976 9469 3985 9503
rect 3985 9469 4019 9503
rect 4019 9469 4028 9503
rect 3976 9460 4028 9469
rect 6920 9571 6972 9580
rect 6920 9537 6929 9571
rect 6929 9537 6963 9571
rect 6963 9537 6972 9571
rect 6920 9528 6972 9537
rect 9312 9528 9364 9580
rect 12164 9571 12216 9580
rect 12164 9537 12173 9571
rect 12173 9537 12207 9571
rect 12207 9537 12216 9571
rect 12164 9528 12216 9537
rect 9036 9503 9088 9512
rect 9036 9469 9045 9503
rect 9045 9469 9079 9503
rect 9079 9469 9088 9503
rect 9036 9460 9088 9469
rect 5356 9392 5408 9444
rect 9956 9392 10008 9444
rect 5264 9324 5316 9376
rect 11428 9324 11480 9376
rect 2514 9222 2566 9274
rect 2578 9222 2630 9274
rect 2642 9222 2694 9274
rect 2706 9222 2758 9274
rect 2770 9222 2822 9274
rect 5642 9222 5694 9274
rect 5706 9222 5758 9274
rect 5770 9222 5822 9274
rect 5834 9222 5886 9274
rect 5898 9222 5950 9274
rect 8770 9222 8822 9274
rect 8834 9222 8886 9274
rect 8898 9222 8950 9274
rect 8962 9222 9014 9274
rect 9026 9222 9078 9274
rect 11898 9222 11950 9274
rect 11962 9222 12014 9274
rect 12026 9222 12078 9274
rect 12090 9222 12142 9274
rect 12154 9222 12206 9274
rect 1768 9120 1820 9172
rect 6276 9120 6328 9172
rect 12440 9120 12492 9172
rect 5264 9027 5316 9036
rect 5264 8993 5273 9027
rect 5273 8993 5307 9027
rect 5307 8993 5316 9027
rect 5264 8984 5316 8993
rect 11428 9027 11480 9036
rect 11428 8993 11437 9027
rect 11437 8993 11471 9027
rect 11471 8993 11480 9027
rect 11428 8984 11480 8993
rect 3056 8959 3108 8968
rect 3056 8925 3065 8959
rect 3065 8925 3099 8959
rect 3099 8925 3108 8959
rect 3056 8916 3108 8925
rect 3240 8959 3292 8968
rect 3240 8925 3249 8959
rect 3249 8925 3283 8959
rect 3283 8925 3292 8959
rect 3240 8916 3292 8925
rect 4988 8959 5040 8968
rect 4988 8925 4997 8959
rect 4997 8925 5031 8959
rect 5031 8925 5040 8959
rect 4988 8916 5040 8925
rect 9496 8916 9548 8968
rect 10232 8916 10284 8968
rect 4620 8848 4672 8900
rect 6920 8848 6972 8900
rect 7564 8848 7616 8900
rect 4712 8780 4764 8832
rect 5356 8780 5408 8832
rect 12716 8848 12768 8900
rect 12900 8780 12952 8832
rect 4078 8678 4130 8730
rect 4142 8678 4194 8730
rect 4206 8678 4258 8730
rect 4270 8678 4322 8730
rect 4334 8678 4386 8730
rect 7206 8678 7258 8730
rect 7270 8678 7322 8730
rect 7334 8678 7386 8730
rect 7398 8678 7450 8730
rect 7462 8678 7514 8730
rect 10334 8678 10386 8730
rect 10398 8678 10450 8730
rect 10462 8678 10514 8730
rect 10526 8678 10578 8730
rect 10590 8678 10642 8730
rect 4988 8576 5040 8628
rect 9496 8576 9548 8628
rect 12808 8619 12860 8628
rect 12808 8585 12817 8619
rect 12817 8585 12851 8619
rect 12851 8585 12860 8619
rect 12808 8576 12860 8585
rect 3976 8483 4028 8492
rect 3976 8449 3985 8483
rect 3985 8449 4019 8483
rect 4019 8449 4028 8483
rect 3976 8440 4028 8449
rect 9128 8440 9180 8492
rect 12624 8483 12676 8492
rect 12624 8449 12633 8483
rect 12633 8449 12667 8483
rect 12667 8449 12676 8483
rect 12624 8440 12676 8449
rect 2514 8134 2566 8186
rect 2578 8134 2630 8186
rect 2642 8134 2694 8186
rect 2706 8134 2758 8186
rect 2770 8134 2822 8186
rect 5642 8134 5694 8186
rect 5706 8134 5758 8186
rect 5770 8134 5822 8186
rect 5834 8134 5886 8186
rect 5898 8134 5950 8186
rect 8770 8134 8822 8186
rect 8834 8134 8886 8186
rect 8898 8134 8950 8186
rect 8962 8134 9014 8186
rect 9026 8134 9078 8186
rect 11898 8134 11950 8186
rect 11962 8134 12014 8186
rect 12026 8134 12078 8186
rect 12090 8134 12142 8186
rect 12154 8134 12206 8186
rect 7012 7896 7064 7948
rect 2044 7828 2096 7880
rect 2320 7871 2372 7880
rect 2320 7837 2329 7871
rect 2329 7837 2363 7871
rect 2363 7837 2372 7871
rect 2320 7828 2372 7837
rect 3976 7828 4028 7880
rect 6920 7828 6972 7880
rect 7656 7828 7708 7880
rect 8300 7828 8352 7880
rect 12900 7939 12952 7948
rect 12900 7905 12909 7939
rect 12909 7905 12943 7939
rect 12943 7905 12952 7939
rect 12900 7896 12952 7905
rect 8944 7871 8996 7880
rect 8944 7837 8953 7871
rect 8953 7837 8987 7871
rect 8987 7837 8996 7871
rect 8944 7828 8996 7837
rect 9496 7760 9548 7812
rect 1492 7735 1544 7744
rect 1492 7701 1501 7735
rect 1501 7701 1535 7735
rect 1535 7701 1544 7735
rect 1492 7692 1544 7701
rect 1676 7692 1728 7744
rect 4436 7692 4488 7744
rect 6644 7735 6696 7744
rect 6644 7701 6653 7735
rect 6653 7701 6687 7735
rect 6687 7701 6696 7735
rect 6644 7692 6696 7701
rect 7104 7692 7156 7744
rect 9588 7692 9640 7744
rect 10692 7735 10744 7744
rect 10692 7701 10701 7735
rect 10701 7701 10735 7735
rect 10735 7701 10744 7735
rect 10692 7692 10744 7701
rect 12348 7760 12400 7812
rect 12808 7692 12860 7744
rect 4078 7590 4130 7642
rect 4142 7590 4194 7642
rect 4206 7590 4258 7642
rect 4270 7590 4322 7642
rect 4334 7590 4386 7642
rect 7206 7590 7258 7642
rect 7270 7590 7322 7642
rect 7334 7590 7386 7642
rect 7398 7590 7450 7642
rect 7462 7590 7514 7642
rect 10334 7590 10386 7642
rect 10398 7590 10450 7642
rect 10462 7590 10514 7642
rect 10526 7590 10578 7642
rect 10590 7590 10642 7642
rect 2044 7488 2096 7540
rect 7564 7488 7616 7540
rect 9496 7488 9548 7540
rect 10968 7531 11020 7540
rect 10968 7497 10977 7531
rect 10977 7497 11011 7531
rect 11011 7497 11020 7531
rect 10968 7488 11020 7497
rect 12716 7531 12768 7540
rect 12716 7497 12725 7531
rect 12725 7497 12759 7531
rect 12759 7497 12768 7531
rect 12716 7488 12768 7497
rect 1676 7463 1728 7472
rect 1676 7429 1685 7463
rect 1685 7429 1719 7463
rect 1719 7429 1728 7463
rect 1676 7420 1728 7429
rect 3884 7420 3936 7472
rect 6644 7463 6696 7472
rect 6644 7429 6653 7463
rect 6653 7429 6687 7463
rect 6687 7429 6696 7463
rect 6644 7420 6696 7429
rect 7104 7420 7156 7472
rect 9588 7420 9640 7472
rect 3608 7395 3660 7404
rect 3608 7361 3617 7395
rect 3617 7361 3651 7395
rect 3651 7361 3660 7395
rect 3608 7352 3660 7361
rect 3976 7352 4028 7404
rect 4436 7395 4488 7404
rect 4436 7361 4445 7395
rect 4445 7361 4479 7395
rect 4479 7361 4488 7395
rect 4436 7352 4488 7361
rect 4896 7352 4948 7404
rect 8300 7352 8352 7404
rect 12808 7395 12860 7404
rect 12808 7361 12817 7395
rect 12817 7361 12851 7395
rect 12851 7361 12860 7395
rect 12808 7352 12860 7361
rect 1400 7327 1452 7336
rect 1400 7293 1409 7327
rect 1409 7293 1443 7327
rect 1443 7293 1452 7327
rect 1400 7284 1452 7293
rect 8944 7284 8996 7336
rect 9864 7284 9916 7336
rect 10692 7284 10744 7336
rect 7012 7148 7064 7200
rect 9588 7148 9640 7200
rect 2514 7046 2566 7098
rect 2578 7046 2630 7098
rect 2642 7046 2694 7098
rect 2706 7046 2758 7098
rect 2770 7046 2822 7098
rect 5642 7046 5694 7098
rect 5706 7046 5758 7098
rect 5770 7046 5822 7098
rect 5834 7046 5886 7098
rect 5898 7046 5950 7098
rect 8770 7046 8822 7098
rect 8834 7046 8886 7098
rect 8898 7046 8950 7098
rect 8962 7046 9014 7098
rect 9026 7046 9078 7098
rect 11898 7046 11950 7098
rect 11962 7046 12014 7098
rect 12026 7046 12078 7098
rect 12090 7046 12142 7098
rect 12154 7046 12206 7098
rect 2320 6987 2372 6996
rect 2320 6953 2329 6987
rect 2329 6953 2363 6987
rect 2363 6953 2372 6987
rect 2320 6944 2372 6953
rect 3976 6944 4028 6996
rect 6920 6987 6972 6996
rect 6920 6953 6929 6987
rect 6929 6953 6963 6987
rect 6963 6953 6972 6987
rect 6920 6944 6972 6953
rect 2412 6808 2464 6860
rect 4896 6808 4948 6860
rect 5264 6808 5316 6860
rect 7564 6851 7616 6860
rect 2044 6740 2096 6792
rect 7564 6817 7573 6851
rect 7573 6817 7607 6851
rect 7607 6817 7616 6851
rect 7564 6808 7616 6817
rect 9864 6876 9916 6928
rect 10232 6808 10284 6860
rect 10876 6808 10928 6860
rect 12348 6808 12400 6860
rect 8576 6740 8628 6792
rect 9312 6740 9364 6792
rect 3516 6604 3568 6656
rect 3884 6604 3936 6656
rect 8300 6672 8352 6724
rect 12808 6672 12860 6724
rect 5724 6647 5776 6656
rect 5724 6613 5733 6647
rect 5733 6613 5767 6647
rect 5767 6613 5776 6647
rect 5724 6604 5776 6613
rect 7656 6604 7708 6656
rect 4078 6502 4130 6554
rect 4142 6502 4194 6554
rect 4206 6502 4258 6554
rect 4270 6502 4322 6554
rect 4334 6502 4386 6554
rect 7206 6502 7258 6554
rect 7270 6502 7322 6554
rect 7334 6502 7386 6554
rect 7398 6502 7450 6554
rect 7462 6502 7514 6554
rect 10334 6502 10386 6554
rect 10398 6502 10450 6554
rect 10462 6502 10514 6554
rect 10526 6502 10578 6554
rect 10590 6502 10642 6554
rect 4528 6400 4580 6452
rect 4620 6400 4672 6452
rect 5264 6400 5316 6452
rect 5724 6400 5776 6452
rect 3884 6332 3936 6384
rect 4712 6332 4764 6384
rect 4896 6307 4948 6316
rect 4896 6273 4905 6307
rect 4905 6273 4939 6307
rect 4939 6273 4948 6307
rect 4896 6264 4948 6273
rect 4620 6239 4672 6248
rect 4620 6205 4629 6239
rect 4629 6205 4663 6239
rect 4663 6205 4672 6239
rect 4620 6196 4672 6205
rect 5724 6128 5776 6180
rect 8300 6400 8352 6452
rect 7104 6332 7156 6384
rect 12992 6196 13044 6248
rect 7656 6128 7708 6180
rect 3516 6060 3568 6112
rect 5540 6060 5592 6112
rect 2514 5958 2566 6010
rect 2578 5958 2630 6010
rect 2642 5958 2694 6010
rect 2706 5958 2758 6010
rect 2770 5958 2822 6010
rect 5642 5958 5694 6010
rect 5706 5958 5758 6010
rect 5770 5958 5822 6010
rect 5834 5958 5886 6010
rect 5898 5958 5950 6010
rect 8770 5958 8822 6010
rect 8834 5958 8886 6010
rect 8898 5958 8950 6010
rect 8962 5958 9014 6010
rect 9026 5958 9078 6010
rect 11898 5958 11950 6010
rect 11962 5958 12014 6010
rect 12026 5958 12078 6010
rect 12090 5958 12142 6010
rect 12154 5958 12206 6010
rect 12808 5831 12860 5840
rect 12808 5797 12817 5831
rect 12817 5797 12851 5831
rect 12851 5797 12860 5831
rect 12808 5788 12860 5797
rect 4620 5720 4672 5772
rect 5172 5720 5224 5772
rect 9680 5763 9732 5772
rect 9680 5729 9689 5763
rect 9689 5729 9723 5763
rect 9723 5729 9732 5763
rect 9680 5720 9732 5729
rect 9864 5652 9916 5704
rect 4528 5584 4580 5636
rect 3884 5559 3936 5568
rect 3884 5525 3893 5559
rect 3893 5525 3927 5559
rect 3927 5525 3936 5559
rect 3884 5516 3936 5525
rect 4436 5516 4488 5568
rect 4712 5516 4764 5568
rect 7656 5516 7708 5568
rect 11336 5695 11388 5704
rect 11336 5661 11345 5695
rect 11345 5661 11379 5695
rect 11379 5661 11388 5695
rect 11336 5652 11388 5661
rect 12532 5652 12584 5704
rect 12808 5652 12860 5704
rect 12624 5627 12676 5636
rect 12624 5593 12633 5627
rect 12633 5593 12667 5627
rect 12667 5593 12676 5627
rect 12624 5584 12676 5593
rect 11428 5516 11480 5568
rect 4078 5414 4130 5466
rect 4142 5414 4194 5466
rect 4206 5414 4258 5466
rect 4270 5414 4322 5466
rect 4334 5414 4386 5466
rect 7206 5414 7258 5466
rect 7270 5414 7322 5466
rect 7334 5414 7386 5466
rect 7398 5414 7450 5466
rect 7462 5414 7514 5466
rect 10334 5414 10386 5466
rect 10398 5414 10450 5466
rect 10462 5414 10514 5466
rect 10526 5414 10578 5466
rect 10590 5414 10642 5466
rect 3976 5312 4028 5364
rect 3884 5176 3936 5228
rect 5540 5312 5592 5364
rect 4712 5244 4764 5296
rect 5172 5219 5224 5228
rect 5172 5185 5181 5219
rect 5181 5185 5215 5219
rect 5215 5185 5224 5219
rect 5172 5176 5224 5185
rect 8116 5312 8168 5364
rect 9588 5312 9640 5364
rect 11336 5312 11388 5364
rect 7564 5244 7616 5296
rect 9312 5244 9364 5296
rect 9680 5244 9732 5296
rect 8668 5108 8720 5160
rect 9588 5219 9640 5228
rect 9220 5108 9272 5160
rect 9588 5185 9597 5219
rect 9597 5185 9631 5219
rect 9631 5185 9640 5219
rect 9588 5176 9640 5185
rect 10692 5219 10744 5228
rect 10692 5185 10701 5219
rect 10701 5185 10735 5219
rect 10735 5185 10744 5219
rect 12624 5219 12676 5228
rect 10692 5176 10744 5185
rect 12624 5185 12633 5219
rect 12633 5185 12667 5219
rect 12667 5185 12676 5219
rect 12624 5176 12676 5185
rect 12716 5108 12768 5160
rect 10784 4972 10836 5024
rect 2514 4870 2566 4922
rect 2578 4870 2630 4922
rect 2642 4870 2694 4922
rect 2706 4870 2758 4922
rect 2770 4870 2822 4922
rect 5642 4870 5694 4922
rect 5706 4870 5758 4922
rect 5770 4870 5822 4922
rect 5834 4870 5886 4922
rect 5898 4870 5950 4922
rect 8770 4870 8822 4922
rect 8834 4870 8886 4922
rect 8898 4870 8950 4922
rect 8962 4870 9014 4922
rect 9026 4870 9078 4922
rect 11898 4870 11950 4922
rect 11962 4870 12014 4922
rect 12026 4870 12078 4922
rect 12090 4870 12142 4922
rect 12154 4870 12206 4922
rect 2136 4607 2188 4616
rect 2136 4573 2145 4607
rect 2145 4573 2179 4607
rect 2179 4573 2188 4607
rect 2136 4564 2188 4573
rect 3240 4564 3292 4616
rect 8668 4632 8720 4684
rect 9220 4675 9272 4684
rect 9220 4641 9229 4675
rect 9229 4641 9263 4675
rect 9263 4641 9272 4675
rect 9220 4632 9272 4641
rect 11428 4675 11480 4684
rect 11428 4641 11437 4675
rect 11437 4641 11471 4675
rect 11471 4641 11480 4675
rect 11428 4632 11480 4641
rect 10232 4564 10284 4616
rect 10692 4564 10744 4616
rect 11152 4607 11204 4616
rect 11152 4573 11161 4607
rect 11161 4573 11195 4607
rect 11195 4573 11204 4607
rect 11152 4564 11204 4573
rect 5448 4496 5500 4548
rect 9220 4496 9272 4548
rect 12716 4496 12768 4548
rect 2872 4428 2924 4480
rect 3792 4428 3844 4480
rect 4712 4471 4764 4480
rect 4712 4437 4721 4471
rect 4721 4437 4755 4471
rect 4755 4437 4764 4471
rect 4712 4428 4764 4437
rect 10692 4471 10744 4480
rect 10692 4437 10701 4471
rect 10701 4437 10735 4471
rect 10735 4437 10744 4471
rect 10692 4428 10744 4437
rect 12808 4428 12860 4480
rect 4078 4326 4130 4378
rect 4142 4326 4194 4378
rect 4206 4326 4258 4378
rect 4270 4326 4322 4378
rect 4334 4326 4386 4378
rect 7206 4326 7258 4378
rect 7270 4326 7322 4378
rect 7334 4326 7386 4378
rect 7398 4326 7450 4378
rect 7462 4326 7514 4378
rect 10334 4326 10386 4378
rect 10398 4326 10450 4378
rect 10462 4326 10514 4378
rect 10526 4326 10578 4378
rect 10590 4326 10642 4378
rect 2136 4224 2188 4276
rect 5172 4224 5224 4276
rect 9220 4267 9272 4276
rect 9220 4233 9229 4267
rect 9229 4233 9263 4267
rect 9263 4233 9272 4267
rect 9220 4224 9272 4233
rect 5448 4156 5500 4208
rect 7564 4156 7616 4208
rect 8668 4156 8720 4208
rect 10232 4156 10284 4208
rect 10692 4199 10744 4208
rect 10692 4165 10701 4199
rect 10701 4165 10735 4199
rect 10735 4165 10744 4199
rect 10692 4156 10744 4165
rect 11152 4224 11204 4276
rect 12716 4267 12768 4276
rect 12716 4233 12725 4267
rect 12725 4233 12759 4267
rect 12759 4233 12768 4267
rect 12716 4224 12768 4233
rect 2320 4131 2372 4140
rect 2320 4097 2329 4131
rect 2329 4097 2363 4131
rect 2363 4097 2372 4131
rect 2320 4088 2372 4097
rect 3240 4131 3292 4140
rect 3240 4097 3249 4131
rect 3249 4097 3283 4131
rect 3283 4097 3292 4131
rect 3240 4088 3292 4097
rect 7012 4131 7064 4140
rect 7012 4097 7021 4131
rect 7021 4097 7055 4131
rect 7055 4097 7064 4131
rect 8116 4131 8168 4140
rect 7012 4088 7064 4097
rect 8116 4097 8125 4131
rect 8125 4097 8159 4131
rect 8159 4097 8168 4131
rect 8116 4088 8168 4097
rect 8576 4131 8628 4140
rect 3148 4020 3200 4072
rect 3516 4063 3568 4072
rect 3516 4029 3525 4063
rect 3525 4029 3559 4063
rect 3559 4029 3568 4063
rect 3516 4020 3568 4029
rect 8576 4097 8585 4131
rect 8585 4097 8619 4131
rect 8619 4097 8628 4131
rect 8576 4088 8628 4097
rect 12900 4131 12952 4140
rect 12900 4097 12909 4131
rect 12909 4097 12943 4131
rect 12943 4097 12952 4131
rect 12900 4088 12952 4097
rect 10692 4020 10744 4072
rect 2412 3884 2464 3936
rect 6552 3927 6604 3936
rect 6552 3893 6561 3927
rect 6561 3893 6595 3927
rect 6595 3893 6604 3927
rect 6552 3884 6604 3893
rect 8668 3884 8720 3936
rect 2514 3782 2566 3834
rect 2578 3782 2630 3834
rect 2642 3782 2694 3834
rect 2706 3782 2758 3834
rect 2770 3782 2822 3834
rect 5642 3782 5694 3834
rect 5706 3782 5758 3834
rect 5770 3782 5822 3834
rect 5834 3782 5886 3834
rect 5898 3782 5950 3834
rect 8770 3782 8822 3834
rect 8834 3782 8886 3834
rect 8898 3782 8950 3834
rect 8962 3782 9014 3834
rect 9026 3782 9078 3834
rect 11898 3782 11950 3834
rect 11962 3782 12014 3834
rect 12026 3782 12078 3834
rect 12090 3782 12142 3834
rect 12154 3782 12206 3834
rect 1676 3680 1728 3732
rect 2320 3680 2372 3732
rect 3608 3680 3660 3732
rect 7564 3723 7616 3732
rect 7564 3689 7573 3723
rect 7573 3689 7607 3723
rect 7607 3689 7616 3723
rect 7564 3680 7616 3689
rect 8576 3680 8628 3732
rect 10692 3723 10744 3732
rect 10692 3689 10701 3723
rect 10701 3689 10735 3723
rect 10735 3689 10744 3723
rect 10692 3680 10744 3689
rect 2872 3587 2924 3596
rect 2872 3553 2881 3587
rect 2881 3553 2915 3587
rect 2915 3553 2924 3587
rect 2872 3544 2924 3553
rect 3792 3519 3844 3528
rect 3792 3485 3801 3519
rect 3801 3485 3835 3519
rect 3835 3485 3844 3519
rect 3792 3476 3844 3485
rect 5448 3476 5500 3528
rect 8668 3544 8720 3596
rect 3424 3408 3476 3460
rect 6368 3408 6420 3460
rect 7104 3340 7156 3392
rect 10784 3408 10836 3460
rect 4078 3238 4130 3290
rect 4142 3238 4194 3290
rect 4206 3238 4258 3290
rect 4270 3238 4322 3290
rect 4334 3238 4386 3290
rect 7206 3238 7258 3290
rect 7270 3238 7322 3290
rect 7334 3238 7386 3290
rect 7398 3238 7450 3290
rect 7462 3238 7514 3290
rect 10334 3238 10386 3290
rect 10398 3238 10450 3290
rect 10462 3238 10514 3290
rect 10526 3238 10578 3290
rect 10590 3238 10642 3290
rect 1492 3179 1544 3188
rect 1492 3145 1501 3179
rect 1501 3145 1535 3179
rect 1535 3145 1544 3179
rect 1492 3136 1544 3145
rect 3516 3136 3568 3188
rect 6368 3179 6420 3188
rect 3424 3068 3476 3120
rect 6368 3145 6377 3179
rect 6377 3145 6411 3179
rect 6411 3145 6420 3179
rect 6368 3136 6420 3145
rect 3792 3068 3844 3120
rect 1676 3043 1728 3052
rect 1676 3009 1685 3043
rect 1685 3009 1719 3043
rect 1719 3009 1728 3043
rect 1676 3000 1728 3009
rect 5356 3068 5408 3120
rect 7104 3068 7156 3120
rect 6552 3043 6604 3052
rect 6552 3009 6561 3043
rect 6561 3009 6595 3043
rect 6595 3009 6604 3043
rect 6552 3000 6604 3009
rect 4712 2932 4764 2984
rect 2514 2694 2566 2746
rect 2578 2694 2630 2746
rect 2642 2694 2694 2746
rect 2706 2694 2758 2746
rect 2770 2694 2822 2746
rect 5642 2694 5694 2746
rect 5706 2694 5758 2746
rect 5770 2694 5822 2746
rect 5834 2694 5886 2746
rect 5898 2694 5950 2746
rect 8770 2694 8822 2746
rect 8834 2694 8886 2746
rect 8898 2694 8950 2746
rect 8962 2694 9014 2746
rect 9026 2694 9078 2746
rect 11898 2694 11950 2746
rect 11962 2694 12014 2746
rect 12026 2694 12078 2746
rect 12090 2694 12142 2746
rect 12154 2694 12206 2746
rect 5448 2592 5500 2644
rect 4436 2524 4488 2576
rect 3240 2456 3292 2508
rect 3884 2388 3936 2440
rect 7564 2388 7616 2440
rect 10692 2388 10744 2440
rect 12808 2388 12860 2440
rect 20 2320 72 2372
rect 7748 2252 7800 2304
rect 11612 2252 11664 2304
rect 12348 2252 12400 2304
rect 4078 2150 4130 2202
rect 4142 2150 4194 2202
rect 4206 2150 4258 2202
rect 4270 2150 4322 2202
rect 4334 2150 4386 2202
rect 7206 2150 7258 2202
rect 7270 2150 7322 2202
rect 7334 2150 7386 2202
rect 7398 2150 7450 2202
rect 7462 2150 7514 2202
rect 10334 2150 10386 2202
rect 10398 2150 10450 2202
rect 10462 2150 10514 2202
rect 10526 2150 10578 2202
rect 10590 2150 10642 2202
<< metal2 >>
rect 2594 16088 2650 16888
rect 6458 16088 6514 16888
rect 10322 16088 10378 16888
rect 14186 16088 14242 16888
rect 1490 15736 1546 15745
rect 1490 15671 1546 15680
rect 1504 14618 1532 15671
rect 2608 14906 2636 16088
rect 2424 14878 2636 14906
rect 1492 14612 1544 14618
rect 1492 14554 1544 14560
rect 2424 14414 2452 14878
rect 2514 14716 2822 14736
rect 2514 14714 2520 14716
rect 2576 14714 2600 14716
rect 2656 14714 2680 14716
rect 2736 14714 2760 14716
rect 2816 14714 2822 14716
rect 2576 14662 2578 14714
rect 2758 14662 2760 14714
rect 2514 14660 2520 14662
rect 2576 14660 2600 14662
rect 2656 14660 2680 14662
rect 2736 14660 2760 14662
rect 2816 14660 2822 14662
rect 2514 14640 2822 14660
rect 5642 14716 5950 14736
rect 5642 14714 5648 14716
rect 5704 14714 5728 14716
rect 5784 14714 5808 14716
rect 5864 14714 5888 14716
rect 5944 14714 5950 14716
rect 5704 14662 5706 14714
rect 5886 14662 5888 14714
rect 5642 14660 5648 14662
rect 5704 14660 5728 14662
rect 5784 14660 5808 14662
rect 5864 14660 5888 14662
rect 5944 14660 5950 14662
rect 5642 14640 5950 14660
rect 6472 14618 6500 16088
rect 8770 14716 9078 14736
rect 8770 14714 8776 14716
rect 8832 14714 8856 14716
rect 8912 14714 8936 14716
rect 8992 14714 9016 14716
rect 9072 14714 9078 14716
rect 8832 14662 8834 14714
rect 9014 14662 9016 14714
rect 8770 14660 8776 14662
rect 8832 14660 8856 14662
rect 8912 14660 8936 14662
rect 8992 14660 9016 14662
rect 9072 14660 9078 14662
rect 8770 14640 9078 14660
rect 10336 14618 10364 16088
rect 11898 14716 12206 14736
rect 11898 14714 11904 14716
rect 11960 14714 11984 14716
rect 12040 14714 12064 14716
rect 12120 14714 12144 14716
rect 12200 14714 12206 14716
rect 11960 14662 11962 14714
rect 12142 14662 12144 14714
rect 11898 14660 11904 14662
rect 11960 14660 11984 14662
rect 12040 14660 12064 14662
rect 12120 14660 12144 14662
rect 12200 14660 12206 14662
rect 11898 14640 12206 14660
rect 14200 14618 14228 16088
rect 6460 14612 6512 14618
rect 6460 14554 6512 14560
rect 10324 14612 10376 14618
rect 10324 14554 10376 14560
rect 14188 14612 14240 14618
rect 14188 14554 14240 14560
rect 2412 14408 2464 14414
rect 2412 14350 2464 14356
rect 7012 14408 7064 14414
rect 7012 14350 7064 14356
rect 10692 14408 10744 14414
rect 10692 14350 10744 14356
rect 12440 14408 12492 14414
rect 12440 14350 12492 14356
rect 3240 14340 3292 14346
rect 3240 14282 3292 14288
rect 2514 13628 2822 13648
rect 2514 13626 2520 13628
rect 2576 13626 2600 13628
rect 2656 13626 2680 13628
rect 2736 13626 2760 13628
rect 2816 13626 2822 13628
rect 2576 13574 2578 13626
rect 2758 13574 2760 13626
rect 2514 13572 2520 13574
rect 2576 13572 2600 13574
rect 2656 13572 2680 13574
rect 2736 13572 2760 13574
rect 2816 13572 2822 13574
rect 2514 13552 2822 13572
rect 2514 12540 2822 12560
rect 2514 12538 2520 12540
rect 2576 12538 2600 12540
rect 2656 12538 2680 12540
rect 2736 12538 2760 12540
rect 2816 12538 2822 12540
rect 2576 12486 2578 12538
rect 2758 12486 2760 12538
rect 2514 12484 2520 12486
rect 2576 12484 2600 12486
rect 2656 12484 2680 12486
rect 2736 12484 2760 12486
rect 2816 12484 2822 12486
rect 2514 12464 2822 12484
rect 2412 11824 2464 11830
rect 2964 11824 3016 11830
rect 2412 11766 2464 11772
rect 2884 11772 2964 11778
rect 2884 11766 3016 11772
rect 2044 11756 2096 11762
rect 2044 11698 2096 11704
rect 1490 11656 1546 11665
rect 1490 11591 1492 11600
rect 1544 11591 1546 11600
rect 1492 11562 1544 11568
rect 2056 11082 2084 11698
rect 2320 11688 2372 11694
rect 2320 11630 2372 11636
rect 2044 11076 2096 11082
rect 2044 11018 2096 11024
rect 2056 10810 2084 11018
rect 2044 10804 2096 10810
rect 2044 10746 2096 10752
rect 2332 10606 2360 11630
rect 2424 11558 2452 11766
rect 2884 11750 3004 11766
rect 2412 11552 2464 11558
rect 2412 11494 2464 11500
rect 1400 10600 1452 10606
rect 1400 10542 1452 10548
rect 2320 10600 2372 10606
rect 2320 10542 2372 10548
rect 1412 9518 1440 10542
rect 1400 9512 1452 9518
rect 1400 9454 1452 9460
rect 1768 9512 1820 9518
rect 1768 9454 1820 9460
rect 1412 7342 1440 9454
rect 1780 9178 1808 9454
rect 1768 9172 1820 9178
rect 1768 9114 1820 9120
rect 2044 7880 2096 7886
rect 2044 7822 2096 7828
rect 2320 7880 2372 7886
rect 2320 7822 2372 7828
rect 1492 7744 1544 7750
rect 1492 7686 1544 7692
rect 1676 7744 1728 7750
rect 1676 7686 1728 7692
rect 1504 7585 1532 7686
rect 1490 7576 1546 7585
rect 1490 7511 1546 7520
rect 1688 7478 1716 7686
rect 2056 7546 2084 7822
rect 2044 7540 2096 7546
rect 2044 7482 2096 7488
rect 1676 7472 1728 7478
rect 1676 7414 1728 7420
rect 1400 7336 1452 7342
rect 1400 7278 1452 7284
rect 2056 6798 2084 7482
rect 2332 7002 2360 7822
rect 2320 6996 2372 7002
rect 2320 6938 2372 6944
rect 2424 6866 2452 11494
rect 2514 11452 2822 11472
rect 2514 11450 2520 11452
rect 2576 11450 2600 11452
rect 2656 11450 2680 11452
rect 2736 11450 2760 11452
rect 2816 11450 2822 11452
rect 2576 11398 2578 11450
rect 2758 11398 2760 11450
rect 2514 11396 2520 11398
rect 2576 11396 2600 11398
rect 2656 11396 2680 11398
rect 2736 11396 2760 11398
rect 2816 11396 2822 11398
rect 2514 11376 2822 11396
rect 2884 10742 2912 11750
rect 2872 10736 2924 10742
rect 2872 10678 2924 10684
rect 2514 10364 2822 10384
rect 2514 10362 2520 10364
rect 2576 10362 2600 10364
rect 2656 10362 2680 10364
rect 2736 10362 2760 10364
rect 2816 10362 2822 10364
rect 2576 10310 2578 10362
rect 2758 10310 2760 10362
rect 2514 10308 2520 10310
rect 2576 10308 2600 10310
rect 2656 10308 2680 10310
rect 2736 10308 2760 10310
rect 2816 10308 2822 10310
rect 2514 10288 2822 10308
rect 2884 9586 2912 10678
rect 3056 9920 3108 9926
rect 3056 9862 3108 9868
rect 2872 9580 2924 9586
rect 2872 9522 2924 9528
rect 2514 9276 2822 9296
rect 2514 9274 2520 9276
rect 2576 9274 2600 9276
rect 2656 9274 2680 9276
rect 2736 9274 2760 9276
rect 2816 9274 2822 9276
rect 2576 9222 2578 9274
rect 2758 9222 2760 9274
rect 2514 9220 2520 9222
rect 2576 9220 2600 9222
rect 2656 9220 2680 9222
rect 2736 9220 2760 9222
rect 2816 9220 2822 9222
rect 2514 9200 2822 9220
rect 3068 8974 3096 9862
rect 3252 9518 3280 14282
rect 4988 14272 5040 14278
rect 4988 14214 5040 14220
rect 4078 14172 4386 14192
rect 4078 14170 4084 14172
rect 4140 14170 4164 14172
rect 4220 14170 4244 14172
rect 4300 14170 4324 14172
rect 4380 14170 4386 14172
rect 4140 14118 4142 14170
rect 4322 14118 4324 14170
rect 4078 14116 4084 14118
rect 4140 14116 4164 14118
rect 4220 14116 4244 14118
rect 4300 14116 4324 14118
rect 4380 14116 4386 14118
rect 4078 14096 4386 14116
rect 4252 13728 4304 13734
rect 4252 13670 4304 13676
rect 4264 13394 4292 13670
rect 4252 13388 4304 13394
rect 4252 13330 4304 13336
rect 4344 13320 4396 13326
rect 4396 13268 4476 13274
rect 4344 13262 4476 13268
rect 4356 13246 4476 13262
rect 4078 13084 4386 13104
rect 4078 13082 4084 13084
rect 4140 13082 4164 13084
rect 4220 13082 4244 13084
rect 4300 13082 4324 13084
rect 4380 13082 4386 13084
rect 4140 13030 4142 13082
rect 4322 13030 4324 13082
rect 4078 13028 4084 13030
rect 4140 13028 4164 13030
rect 4220 13028 4244 13030
rect 4300 13028 4324 13030
rect 4380 13028 4386 13030
rect 4078 13008 4386 13028
rect 4448 12306 4476 13246
rect 5000 12850 5028 14214
rect 6368 13932 6420 13938
rect 6368 13874 6420 13880
rect 5642 13628 5950 13648
rect 5642 13626 5648 13628
rect 5704 13626 5728 13628
rect 5784 13626 5808 13628
rect 5864 13626 5888 13628
rect 5944 13626 5950 13628
rect 5704 13574 5706 13626
rect 5886 13574 5888 13626
rect 5642 13572 5648 13574
rect 5704 13572 5728 13574
rect 5784 13572 5808 13574
rect 5864 13572 5888 13574
rect 5944 13572 5950 13574
rect 5642 13552 5950 13572
rect 5448 13184 5500 13190
rect 5448 13126 5500 13132
rect 5460 12850 5488 13126
rect 6380 12986 6408 13874
rect 6828 13728 6880 13734
rect 6828 13670 6880 13676
rect 6840 13394 6868 13670
rect 6828 13388 6880 13394
rect 6828 13330 6880 13336
rect 6552 13320 6604 13326
rect 6552 13262 6604 13268
rect 6368 12980 6420 12986
rect 6368 12922 6420 12928
rect 4988 12844 5040 12850
rect 4988 12786 5040 12792
rect 5264 12844 5316 12850
rect 5264 12786 5316 12792
rect 5448 12844 5500 12850
rect 5448 12786 5500 12792
rect 4896 12640 4948 12646
rect 4896 12582 4948 12588
rect 4908 12306 4936 12582
rect 4436 12300 4488 12306
rect 4436 12242 4488 12248
rect 4620 12300 4672 12306
rect 4620 12242 4672 12248
rect 4896 12300 4948 12306
rect 4896 12242 4948 12248
rect 4078 11996 4386 12016
rect 4078 11994 4084 11996
rect 4140 11994 4164 11996
rect 4220 11994 4244 11996
rect 4300 11994 4324 11996
rect 4380 11994 4386 11996
rect 4140 11942 4142 11994
rect 4322 11942 4324 11994
rect 4078 11940 4084 11942
rect 4140 11940 4164 11942
rect 4220 11940 4244 11942
rect 4300 11940 4324 11942
rect 4380 11940 4386 11942
rect 4078 11920 4386 11940
rect 4160 11688 4212 11694
rect 4160 11630 4212 11636
rect 4172 11150 4200 11630
rect 4160 11144 4212 11150
rect 4160 11086 4212 11092
rect 4436 11144 4488 11150
rect 4436 11086 4488 11092
rect 3792 11008 3844 11014
rect 3792 10950 3844 10956
rect 3804 10742 3832 10950
rect 4078 10908 4386 10928
rect 4078 10906 4084 10908
rect 4140 10906 4164 10908
rect 4220 10906 4244 10908
rect 4300 10906 4324 10908
rect 4380 10906 4386 10908
rect 4140 10854 4142 10906
rect 4322 10854 4324 10906
rect 4078 10852 4084 10854
rect 4140 10852 4164 10854
rect 4220 10852 4244 10854
rect 4300 10852 4324 10854
rect 4380 10852 4386 10854
rect 4078 10832 4386 10852
rect 3792 10736 3844 10742
rect 3792 10678 3844 10684
rect 4448 10130 4476 11086
rect 4436 10124 4488 10130
rect 4436 10066 4488 10072
rect 4632 10062 4660 12242
rect 5276 11694 5304 12786
rect 6276 12708 6328 12714
rect 6276 12650 6328 12656
rect 5642 12540 5950 12560
rect 5642 12538 5648 12540
rect 5704 12538 5728 12540
rect 5784 12538 5808 12540
rect 5864 12538 5888 12540
rect 5944 12538 5950 12540
rect 5704 12486 5706 12538
rect 5886 12486 5888 12538
rect 5642 12484 5648 12486
rect 5704 12484 5728 12486
rect 5784 12484 5808 12486
rect 5864 12484 5888 12486
rect 5944 12484 5950 12486
rect 5642 12464 5950 12484
rect 6288 12442 6316 12650
rect 6276 12436 6328 12442
rect 6276 12378 6328 12384
rect 6564 11762 6592 13262
rect 6552 11756 6604 11762
rect 6552 11698 6604 11704
rect 5264 11688 5316 11694
rect 5264 11630 5316 11636
rect 5642 11452 5950 11472
rect 5642 11450 5648 11452
rect 5704 11450 5728 11452
rect 5784 11450 5808 11452
rect 5864 11450 5888 11452
rect 5944 11450 5950 11452
rect 5704 11398 5706 11450
rect 5886 11398 5888 11450
rect 5642 11396 5648 11398
rect 5704 11396 5728 11398
rect 5784 11396 5808 11398
rect 5864 11396 5888 11398
rect 5944 11396 5950 11398
rect 5642 11376 5950 11396
rect 6564 11218 6592 11698
rect 6552 11212 6604 11218
rect 6552 11154 6604 11160
rect 5642 10364 5950 10384
rect 5642 10362 5648 10364
rect 5704 10362 5728 10364
rect 5784 10362 5808 10364
rect 5864 10362 5888 10364
rect 5944 10362 5950 10364
rect 5704 10310 5706 10362
rect 5886 10310 5888 10362
rect 5642 10308 5648 10310
rect 5704 10308 5728 10310
rect 5784 10308 5808 10310
rect 5864 10308 5888 10310
rect 5944 10308 5950 10310
rect 5642 10288 5950 10308
rect 6276 10260 6328 10266
rect 6276 10202 6328 10208
rect 4620 10056 4672 10062
rect 4620 9998 4672 10004
rect 4988 10056 5040 10062
rect 4988 9998 5040 10004
rect 4528 9920 4580 9926
rect 4528 9862 4580 9868
rect 4078 9820 4386 9840
rect 4078 9818 4084 9820
rect 4140 9818 4164 9820
rect 4220 9818 4244 9820
rect 4300 9818 4324 9820
rect 4380 9818 4386 9820
rect 4140 9766 4142 9818
rect 4322 9766 4324 9818
rect 4078 9764 4084 9766
rect 4140 9764 4164 9766
rect 4220 9764 4244 9766
rect 4300 9764 4324 9766
rect 4380 9764 4386 9766
rect 4078 9744 4386 9764
rect 4540 9654 4568 9862
rect 4528 9648 4580 9654
rect 4528 9590 4580 9596
rect 3240 9512 3292 9518
rect 3240 9454 3292 9460
rect 3976 9512 4028 9518
rect 3976 9454 4028 9460
rect 3252 8974 3280 9454
rect 3056 8968 3108 8974
rect 3056 8910 3108 8916
rect 3240 8968 3292 8974
rect 3240 8910 3292 8916
rect 2514 8188 2822 8208
rect 2514 8186 2520 8188
rect 2576 8186 2600 8188
rect 2656 8186 2680 8188
rect 2736 8186 2760 8188
rect 2816 8186 2822 8188
rect 2576 8134 2578 8186
rect 2758 8134 2760 8186
rect 2514 8132 2520 8134
rect 2576 8132 2600 8134
rect 2656 8132 2680 8134
rect 2736 8132 2760 8134
rect 2816 8132 2822 8134
rect 2514 8112 2822 8132
rect 2514 7100 2822 7120
rect 2514 7098 2520 7100
rect 2576 7098 2600 7100
rect 2656 7098 2680 7100
rect 2736 7098 2760 7100
rect 2816 7098 2822 7100
rect 2576 7046 2578 7098
rect 2758 7046 2760 7098
rect 2514 7044 2520 7046
rect 2576 7044 2600 7046
rect 2656 7044 2680 7046
rect 2736 7044 2760 7046
rect 2816 7044 2822 7046
rect 2514 7024 2822 7044
rect 3252 6914 3280 8910
rect 3988 8498 4016 9454
rect 4078 8732 4386 8752
rect 4078 8730 4084 8732
rect 4140 8730 4164 8732
rect 4220 8730 4244 8732
rect 4300 8730 4324 8732
rect 4380 8730 4386 8732
rect 4140 8678 4142 8730
rect 4322 8678 4324 8730
rect 4078 8676 4084 8678
rect 4140 8676 4164 8678
rect 4220 8676 4244 8678
rect 4300 8676 4324 8678
rect 4380 8676 4386 8678
rect 4078 8656 4386 8676
rect 3976 8492 4028 8498
rect 3976 8434 4028 8440
rect 3988 7886 4016 8434
rect 3976 7880 4028 7886
rect 3976 7822 4028 7828
rect 3884 7472 3936 7478
rect 3884 7414 3936 7420
rect 3608 7404 3660 7410
rect 3608 7346 3660 7352
rect 3160 6886 3280 6914
rect 2412 6860 2464 6866
rect 2412 6802 2464 6808
rect 2044 6792 2096 6798
rect 2044 6734 2096 6740
rect 2136 4616 2188 4622
rect 2136 4558 2188 4564
rect 2148 4282 2176 4558
rect 2136 4276 2188 4282
rect 2136 4218 2188 4224
rect 2320 4140 2372 4146
rect 2320 4082 2372 4088
rect 2332 3738 2360 4082
rect 2424 3942 2452 6802
rect 2514 6012 2822 6032
rect 2514 6010 2520 6012
rect 2576 6010 2600 6012
rect 2656 6010 2680 6012
rect 2736 6010 2760 6012
rect 2816 6010 2822 6012
rect 2576 5958 2578 6010
rect 2758 5958 2760 6010
rect 2514 5956 2520 5958
rect 2576 5956 2600 5958
rect 2656 5956 2680 5958
rect 2736 5956 2760 5958
rect 2816 5956 2822 5958
rect 2514 5936 2822 5956
rect 2514 4924 2822 4944
rect 2514 4922 2520 4924
rect 2576 4922 2600 4924
rect 2656 4922 2680 4924
rect 2736 4922 2760 4924
rect 2816 4922 2822 4924
rect 2576 4870 2578 4922
rect 2758 4870 2760 4922
rect 2514 4868 2520 4870
rect 2576 4868 2600 4870
rect 2656 4868 2680 4870
rect 2736 4868 2760 4870
rect 2816 4868 2822 4870
rect 2514 4848 2822 4868
rect 2872 4480 2924 4486
rect 2872 4422 2924 4428
rect 2412 3936 2464 3942
rect 2412 3878 2464 3884
rect 2514 3836 2822 3856
rect 2514 3834 2520 3836
rect 2576 3834 2600 3836
rect 2656 3834 2680 3836
rect 2736 3834 2760 3836
rect 2816 3834 2822 3836
rect 2576 3782 2578 3834
rect 2758 3782 2760 3834
rect 2514 3780 2520 3782
rect 2576 3780 2600 3782
rect 2656 3780 2680 3782
rect 2736 3780 2760 3782
rect 2816 3780 2822 3782
rect 2514 3760 2822 3780
rect 1676 3732 1728 3738
rect 1676 3674 1728 3680
rect 2320 3732 2372 3738
rect 2320 3674 2372 3680
rect 1490 3496 1546 3505
rect 1490 3431 1546 3440
rect 1504 3194 1532 3431
rect 1492 3188 1544 3194
rect 1492 3130 1544 3136
rect 1688 3058 1716 3674
rect 2884 3602 2912 4422
rect 3160 4078 3188 6886
rect 3516 6656 3568 6662
rect 3516 6598 3568 6604
rect 3528 6118 3556 6598
rect 3516 6112 3568 6118
rect 3516 6054 3568 6060
rect 3240 4616 3292 4622
rect 3240 4558 3292 4564
rect 3252 4146 3280 4558
rect 3240 4140 3292 4146
rect 3240 4082 3292 4088
rect 3148 4072 3200 4078
rect 3148 4014 3200 4020
rect 2872 3596 2924 3602
rect 2872 3538 2924 3544
rect 1676 3052 1728 3058
rect 1676 2994 1728 3000
rect 2514 2748 2822 2768
rect 2514 2746 2520 2748
rect 2576 2746 2600 2748
rect 2656 2746 2680 2748
rect 2736 2746 2760 2748
rect 2816 2746 2822 2748
rect 2576 2694 2578 2746
rect 2758 2694 2760 2746
rect 2514 2692 2520 2694
rect 2576 2692 2600 2694
rect 2656 2692 2680 2694
rect 2736 2692 2760 2694
rect 2816 2692 2822 2694
rect 2514 2672 2822 2692
rect 3252 2514 3280 4082
rect 3516 4072 3568 4078
rect 3516 4014 3568 4020
rect 3424 3460 3476 3466
rect 3424 3402 3476 3408
rect 3436 3126 3464 3402
rect 3528 3194 3556 4014
rect 3620 3738 3648 7346
rect 3896 6662 3924 7414
rect 3988 7410 4016 7822
rect 4436 7744 4488 7750
rect 4436 7686 4488 7692
rect 4078 7644 4386 7664
rect 4078 7642 4084 7644
rect 4140 7642 4164 7644
rect 4220 7642 4244 7644
rect 4300 7642 4324 7644
rect 4380 7642 4386 7644
rect 4140 7590 4142 7642
rect 4322 7590 4324 7642
rect 4078 7588 4084 7590
rect 4140 7588 4164 7590
rect 4220 7588 4244 7590
rect 4300 7588 4324 7590
rect 4380 7588 4386 7590
rect 4078 7568 4386 7588
rect 4448 7410 4476 7686
rect 3976 7404 4028 7410
rect 3976 7346 4028 7352
rect 4436 7404 4488 7410
rect 4436 7346 4488 7352
rect 3976 6996 4028 7002
rect 3976 6938 4028 6944
rect 3884 6656 3936 6662
rect 3884 6598 3936 6604
rect 3896 6390 3924 6598
rect 3884 6384 3936 6390
rect 3884 6326 3936 6332
rect 3884 5568 3936 5574
rect 3884 5510 3936 5516
rect 3896 5234 3924 5510
rect 3988 5370 4016 6938
rect 4078 6556 4386 6576
rect 4078 6554 4084 6556
rect 4140 6554 4164 6556
rect 4220 6554 4244 6556
rect 4300 6554 4324 6556
rect 4380 6554 4386 6556
rect 4140 6502 4142 6554
rect 4322 6502 4324 6554
rect 4078 6500 4084 6502
rect 4140 6500 4164 6502
rect 4220 6500 4244 6502
rect 4300 6500 4324 6502
rect 4380 6500 4386 6502
rect 4078 6480 4386 6500
rect 4540 6458 4568 9590
rect 5000 8974 5028 9998
rect 6288 9994 6316 10202
rect 6276 9988 6328 9994
rect 6276 9930 6328 9936
rect 5356 9444 5408 9450
rect 5356 9386 5408 9392
rect 5264 9376 5316 9382
rect 5264 9318 5316 9324
rect 5276 9042 5304 9318
rect 5264 9036 5316 9042
rect 5264 8978 5316 8984
rect 4988 8968 5040 8974
rect 4988 8910 5040 8916
rect 4620 8900 4672 8906
rect 4620 8842 4672 8848
rect 4632 6458 4660 8842
rect 4712 8832 4764 8838
rect 4712 8774 4764 8780
rect 4528 6452 4580 6458
rect 4528 6394 4580 6400
rect 4620 6452 4672 6458
rect 4620 6394 4672 6400
rect 4632 6338 4660 6394
rect 4724 6390 4752 8774
rect 5000 8634 5028 8910
rect 5368 8838 5396 9386
rect 5642 9276 5950 9296
rect 5642 9274 5648 9276
rect 5704 9274 5728 9276
rect 5784 9274 5808 9276
rect 5864 9274 5888 9276
rect 5944 9274 5950 9276
rect 5704 9222 5706 9274
rect 5886 9222 5888 9274
rect 5642 9220 5648 9222
rect 5704 9220 5728 9222
rect 5784 9220 5808 9222
rect 5864 9220 5888 9222
rect 5944 9220 5950 9222
rect 5642 9200 5950 9220
rect 6288 9178 6316 9930
rect 6564 9926 6592 11154
rect 6920 11076 6972 11082
rect 6920 11018 6972 11024
rect 6932 10266 6960 11018
rect 6920 10260 6972 10266
rect 6920 10202 6972 10208
rect 6920 9988 6972 9994
rect 6920 9930 6972 9936
rect 6552 9920 6604 9926
rect 6552 9862 6604 9868
rect 6932 9586 6960 9930
rect 6920 9580 6972 9586
rect 6920 9522 6972 9528
rect 6276 9172 6328 9178
rect 6276 9114 6328 9120
rect 6932 8906 6960 9522
rect 6920 8900 6972 8906
rect 6920 8842 6972 8848
rect 5356 8832 5408 8838
rect 5356 8774 5408 8780
rect 4988 8628 5040 8634
rect 4988 8570 5040 8576
rect 5642 8188 5950 8208
rect 5642 8186 5648 8188
rect 5704 8186 5728 8188
rect 5784 8186 5808 8188
rect 5864 8186 5888 8188
rect 5944 8186 5950 8188
rect 5704 8134 5706 8186
rect 5886 8134 5888 8186
rect 5642 8132 5648 8134
rect 5704 8132 5728 8134
rect 5784 8132 5808 8134
rect 5864 8132 5888 8134
rect 5944 8132 5950 8134
rect 5642 8112 5950 8132
rect 7024 7954 7052 14350
rect 7206 14172 7514 14192
rect 7206 14170 7212 14172
rect 7268 14170 7292 14172
rect 7348 14170 7372 14172
rect 7428 14170 7452 14172
rect 7508 14170 7514 14172
rect 7268 14118 7270 14170
rect 7450 14118 7452 14170
rect 7206 14116 7212 14118
rect 7268 14116 7292 14118
rect 7348 14116 7372 14118
rect 7428 14116 7452 14118
rect 7508 14116 7514 14118
rect 7206 14096 7514 14116
rect 10334 14172 10642 14192
rect 10334 14170 10340 14172
rect 10396 14170 10420 14172
rect 10476 14170 10500 14172
rect 10556 14170 10580 14172
rect 10636 14170 10642 14172
rect 10396 14118 10398 14170
rect 10578 14118 10580 14170
rect 10334 14116 10340 14118
rect 10396 14116 10420 14118
rect 10476 14116 10500 14118
rect 10556 14116 10580 14118
rect 10636 14116 10642 14118
rect 10334 14096 10642 14116
rect 9772 13932 9824 13938
rect 9772 13874 9824 13880
rect 10232 13932 10284 13938
rect 10232 13874 10284 13880
rect 9220 13728 9272 13734
rect 9220 13670 9272 13676
rect 8770 13628 9078 13648
rect 8770 13626 8776 13628
rect 8832 13626 8856 13628
rect 8912 13626 8936 13628
rect 8992 13626 9016 13628
rect 9072 13626 9078 13628
rect 8832 13574 8834 13626
rect 9014 13574 9016 13626
rect 8770 13572 8776 13574
rect 8832 13572 8856 13574
rect 8912 13572 8936 13574
rect 8992 13572 9016 13574
rect 9072 13572 9078 13574
rect 8770 13552 9078 13572
rect 9232 13394 9260 13670
rect 9220 13388 9272 13394
rect 9220 13330 9272 13336
rect 8208 13252 8260 13258
rect 8208 13194 8260 13200
rect 7206 13084 7514 13104
rect 7206 13082 7212 13084
rect 7268 13082 7292 13084
rect 7348 13082 7372 13084
rect 7428 13082 7452 13084
rect 7508 13082 7514 13084
rect 7268 13030 7270 13082
rect 7450 13030 7452 13082
rect 7206 13028 7212 13030
rect 7268 13028 7292 13030
rect 7348 13028 7372 13030
rect 7428 13028 7452 13030
rect 7508 13028 7514 13030
rect 7206 13008 7514 13028
rect 8220 12170 8248 13194
rect 8300 13184 8352 13190
rect 8300 13126 8352 13132
rect 9588 13184 9640 13190
rect 9588 13126 9640 13132
rect 8208 12164 8260 12170
rect 8208 12106 8260 12112
rect 7932 12096 7984 12102
rect 7932 12038 7984 12044
rect 7206 11996 7514 12016
rect 7206 11994 7212 11996
rect 7268 11994 7292 11996
rect 7348 11994 7372 11996
rect 7428 11994 7452 11996
rect 7508 11994 7514 11996
rect 7268 11942 7270 11994
rect 7450 11942 7452 11994
rect 7206 11940 7212 11942
rect 7268 11940 7292 11942
rect 7348 11940 7372 11942
rect 7428 11940 7452 11942
rect 7508 11940 7514 11942
rect 7206 11920 7514 11940
rect 7944 11558 7972 12038
rect 7932 11552 7984 11558
rect 7932 11494 7984 11500
rect 8220 11082 8248 12106
rect 8208 11076 8260 11082
rect 8208 11018 8260 11024
rect 7206 10908 7514 10928
rect 7206 10906 7212 10908
rect 7268 10906 7292 10908
rect 7348 10906 7372 10908
rect 7428 10906 7452 10908
rect 7508 10906 7514 10908
rect 7268 10854 7270 10906
rect 7450 10854 7452 10906
rect 7206 10852 7212 10854
rect 7268 10852 7292 10854
rect 7348 10852 7372 10854
rect 7428 10852 7452 10854
rect 7508 10852 7514 10854
rect 7206 10832 7514 10852
rect 8312 10742 8340 13126
rect 8770 12540 9078 12560
rect 8770 12538 8776 12540
rect 8832 12538 8856 12540
rect 8912 12538 8936 12540
rect 8992 12538 9016 12540
rect 9072 12538 9078 12540
rect 8832 12486 8834 12538
rect 9014 12486 9016 12538
rect 8770 12484 8776 12486
rect 8832 12484 8856 12486
rect 8912 12484 8936 12486
rect 8992 12484 9016 12486
rect 9072 12484 9078 12486
rect 8770 12464 9078 12484
rect 9600 12238 9628 13126
rect 9784 12986 9812 13874
rect 10048 13864 10100 13870
rect 10048 13806 10100 13812
rect 9772 12980 9824 12986
rect 9772 12922 9824 12928
rect 9588 12232 9640 12238
rect 9588 12174 9640 12180
rect 9128 12164 9180 12170
rect 9128 12106 9180 12112
rect 9140 11898 9168 12106
rect 9128 11892 9180 11898
rect 9128 11834 9180 11840
rect 8392 11688 8444 11694
rect 8392 11630 8444 11636
rect 8404 11354 8432 11630
rect 8770 11452 9078 11472
rect 8770 11450 8776 11452
rect 8832 11450 8856 11452
rect 8912 11450 8936 11452
rect 8992 11450 9016 11452
rect 9072 11450 9078 11452
rect 8832 11398 8834 11450
rect 9014 11398 9016 11450
rect 8770 11396 8776 11398
rect 8832 11396 8856 11398
rect 8912 11396 8936 11398
rect 8992 11396 9016 11398
rect 9072 11396 9078 11398
rect 8770 11376 9078 11396
rect 8392 11348 8444 11354
rect 8392 11290 8444 11296
rect 8300 10736 8352 10742
rect 8300 10678 8352 10684
rect 7656 10600 7708 10606
rect 7656 10542 7708 10548
rect 7668 10266 7696 10542
rect 8116 10464 8168 10470
rect 8116 10406 8168 10412
rect 7656 10260 7708 10266
rect 7656 10202 7708 10208
rect 8128 10130 8156 10406
rect 8116 10124 8168 10130
rect 8116 10066 8168 10072
rect 7206 9820 7514 9840
rect 7206 9818 7212 9820
rect 7268 9818 7292 9820
rect 7348 9818 7372 9820
rect 7428 9818 7452 9820
rect 7508 9818 7514 9820
rect 7268 9766 7270 9818
rect 7450 9766 7452 9818
rect 7206 9764 7212 9766
rect 7268 9764 7292 9766
rect 7348 9764 7372 9766
rect 7428 9764 7452 9766
rect 7508 9764 7514 9766
rect 7206 9744 7514 9764
rect 7564 8900 7616 8906
rect 7564 8842 7616 8848
rect 7206 8732 7514 8752
rect 7206 8730 7212 8732
rect 7268 8730 7292 8732
rect 7348 8730 7372 8732
rect 7428 8730 7452 8732
rect 7508 8730 7514 8732
rect 7268 8678 7270 8730
rect 7450 8678 7452 8730
rect 7206 8676 7212 8678
rect 7268 8676 7292 8678
rect 7348 8676 7372 8678
rect 7428 8676 7452 8678
rect 7508 8676 7514 8678
rect 7206 8656 7514 8676
rect 7012 7948 7064 7954
rect 7012 7890 7064 7896
rect 6920 7880 6972 7886
rect 6920 7822 6972 7828
rect 6644 7744 6696 7750
rect 6644 7686 6696 7692
rect 6656 7478 6684 7686
rect 6644 7472 6696 7478
rect 6644 7414 6696 7420
rect 4896 7404 4948 7410
rect 4896 7346 4948 7352
rect 4908 6866 4936 7346
rect 5642 7100 5950 7120
rect 5642 7098 5648 7100
rect 5704 7098 5728 7100
rect 5784 7098 5808 7100
rect 5864 7098 5888 7100
rect 5944 7098 5950 7100
rect 5704 7046 5706 7098
rect 5886 7046 5888 7098
rect 5642 7044 5648 7046
rect 5704 7044 5728 7046
rect 5784 7044 5808 7046
rect 5864 7044 5888 7046
rect 5944 7044 5950 7046
rect 5642 7024 5950 7044
rect 6932 7002 6960 7822
rect 7024 7206 7052 7890
rect 7104 7744 7156 7750
rect 7104 7686 7156 7692
rect 7116 7478 7144 7686
rect 7206 7644 7514 7664
rect 7206 7642 7212 7644
rect 7268 7642 7292 7644
rect 7348 7642 7372 7644
rect 7428 7642 7452 7644
rect 7508 7642 7514 7644
rect 7268 7590 7270 7642
rect 7450 7590 7452 7642
rect 7206 7588 7212 7590
rect 7268 7588 7292 7590
rect 7348 7588 7372 7590
rect 7428 7588 7452 7590
rect 7508 7588 7514 7590
rect 7206 7568 7514 7588
rect 7576 7546 7604 8842
rect 7656 7880 7708 7886
rect 7656 7822 7708 7828
rect 7564 7540 7616 7546
rect 7564 7482 7616 7488
rect 7104 7472 7156 7478
rect 7668 7426 7696 7822
rect 7104 7414 7156 7420
rect 7012 7200 7064 7206
rect 7012 7142 7064 7148
rect 6920 6996 6972 7002
rect 6920 6938 6972 6944
rect 4896 6860 4948 6866
rect 4896 6802 4948 6808
rect 5264 6860 5316 6866
rect 5264 6802 5316 6808
rect 4540 6310 4660 6338
rect 4712 6384 4764 6390
rect 4712 6326 4764 6332
rect 4540 5642 4568 6310
rect 4620 6248 4672 6254
rect 4620 6190 4672 6196
rect 4632 5778 4660 6190
rect 4620 5772 4672 5778
rect 4620 5714 4672 5720
rect 4528 5636 4580 5642
rect 4528 5578 4580 5584
rect 4724 5574 4752 6326
rect 4908 6322 4936 6802
rect 5276 6458 5304 6802
rect 5724 6656 5776 6662
rect 5724 6598 5776 6604
rect 5736 6458 5764 6598
rect 5264 6452 5316 6458
rect 5264 6394 5316 6400
rect 5724 6452 5776 6458
rect 5724 6394 5776 6400
rect 4896 6316 4948 6322
rect 4896 6258 4948 6264
rect 5736 6186 5764 6394
rect 5724 6180 5776 6186
rect 5724 6122 5776 6128
rect 5540 6112 5592 6118
rect 5540 6054 5592 6060
rect 5172 5772 5224 5778
rect 5172 5714 5224 5720
rect 4436 5568 4488 5574
rect 4436 5510 4488 5516
rect 4712 5568 4764 5574
rect 4712 5510 4764 5516
rect 4078 5468 4386 5488
rect 4078 5466 4084 5468
rect 4140 5466 4164 5468
rect 4220 5466 4244 5468
rect 4300 5466 4324 5468
rect 4380 5466 4386 5468
rect 4140 5414 4142 5466
rect 4322 5414 4324 5466
rect 4078 5412 4084 5414
rect 4140 5412 4164 5414
rect 4220 5412 4244 5414
rect 4300 5412 4324 5414
rect 4380 5412 4386 5414
rect 4078 5392 4386 5412
rect 3976 5364 4028 5370
rect 3976 5306 4028 5312
rect 3884 5228 3936 5234
rect 3884 5170 3936 5176
rect 3792 4480 3844 4486
rect 3792 4422 3844 4428
rect 3608 3732 3660 3738
rect 3608 3674 3660 3680
rect 3804 3534 3832 4422
rect 4078 4380 4386 4400
rect 4078 4378 4084 4380
rect 4140 4378 4164 4380
rect 4220 4378 4244 4380
rect 4300 4378 4324 4380
rect 4380 4378 4386 4380
rect 4140 4326 4142 4378
rect 4322 4326 4324 4378
rect 4078 4324 4084 4326
rect 4140 4324 4164 4326
rect 4220 4324 4244 4326
rect 4300 4324 4324 4326
rect 4380 4324 4386 4326
rect 4078 4304 4386 4324
rect 3792 3528 3844 3534
rect 3792 3470 3844 3476
rect 3516 3188 3568 3194
rect 3516 3130 3568 3136
rect 3804 3126 3832 3470
rect 4078 3292 4386 3312
rect 4078 3290 4084 3292
rect 4140 3290 4164 3292
rect 4220 3290 4244 3292
rect 4300 3290 4324 3292
rect 4380 3290 4386 3292
rect 4140 3238 4142 3290
rect 4322 3238 4324 3290
rect 4078 3236 4084 3238
rect 4140 3236 4164 3238
rect 4220 3236 4244 3238
rect 4300 3236 4324 3238
rect 4380 3236 4386 3238
rect 4078 3216 4386 3236
rect 3424 3120 3476 3126
rect 3424 3062 3476 3068
rect 3792 3120 3844 3126
rect 3792 3062 3844 3068
rect 4448 2582 4476 5510
rect 4712 5296 4764 5302
rect 4712 5238 4764 5244
rect 4724 4486 4752 5238
rect 5184 5234 5212 5714
rect 5552 5370 5580 6054
rect 5642 6012 5950 6032
rect 5642 6010 5648 6012
rect 5704 6010 5728 6012
rect 5784 6010 5808 6012
rect 5864 6010 5888 6012
rect 5944 6010 5950 6012
rect 5704 5958 5706 6010
rect 5886 5958 5888 6010
rect 5642 5956 5648 5958
rect 5704 5956 5728 5958
rect 5784 5956 5808 5958
rect 5864 5956 5888 5958
rect 5944 5956 5950 5958
rect 5642 5936 5950 5956
rect 5540 5364 5592 5370
rect 5540 5306 5592 5312
rect 5172 5228 5224 5234
rect 5172 5170 5224 5176
rect 4712 4480 4764 4486
rect 4712 4422 4764 4428
rect 4724 2990 4752 4422
rect 5184 4282 5212 5170
rect 5642 4924 5950 4944
rect 5642 4922 5648 4924
rect 5704 4922 5728 4924
rect 5784 4922 5808 4924
rect 5864 4922 5888 4924
rect 5944 4922 5950 4924
rect 5704 4870 5706 4922
rect 5886 4870 5888 4922
rect 5642 4868 5648 4870
rect 5704 4868 5728 4870
rect 5784 4868 5808 4870
rect 5864 4868 5888 4870
rect 5944 4868 5950 4870
rect 5642 4848 5950 4868
rect 5448 4548 5500 4554
rect 5448 4490 5500 4496
rect 5172 4276 5224 4282
rect 5172 4218 5224 4224
rect 5460 4214 5488 4490
rect 5448 4208 5500 4214
rect 5448 4150 5500 4156
rect 5460 3618 5488 4150
rect 7024 4146 7052 7142
rect 7116 6390 7144 7414
rect 7576 7398 7696 7426
rect 7576 6866 7604 7398
rect 7564 6860 7616 6866
rect 7564 6802 7616 6808
rect 7206 6556 7514 6576
rect 7206 6554 7212 6556
rect 7268 6554 7292 6556
rect 7348 6554 7372 6556
rect 7428 6554 7452 6556
rect 7508 6554 7514 6556
rect 7268 6502 7270 6554
rect 7450 6502 7452 6554
rect 7206 6500 7212 6502
rect 7268 6500 7292 6502
rect 7348 6500 7372 6502
rect 7428 6500 7452 6502
rect 7508 6500 7514 6502
rect 7206 6480 7514 6500
rect 7104 6384 7156 6390
rect 7104 6326 7156 6332
rect 7206 5468 7514 5488
rect 7206 5466 7212 5468
rect 7268 5466 7292 5468
rect 7348 5466 7372 5468
rect 7428 5466 7452 5468
rect 7508 5466 7514 5468
rect 7268 5414 7270 5466
rect 7450 5414 7452 5466
rect 7206 5412 7212 5414
rect 7268 5412 7292 5414
rect 7348 5412 7372 5414
rect 7428 5412 7452 5414
rect 7508 5412 7514 5414
rect 7206 5392 7514 5412
rect 7576 5302 7604 6802
rect 7656 6656 7708 6662
rect 7656 6598 7708 6604
rect 7668 6186 7696 6598
rect 7656 6180 7708 6186
rect 7656 6122 7708 6128
rect 7668 5574 7696 6122
rect 7656 5568 7708 5574
rect 7656 5510 7708 5516
rect 8128 5370 8156 10066
rect 8312 7886 8340 10678
rect 9140 10674 9168 11834
rect 9600 11558 9628 12174
rect 10060 12102 10088 13806
rect 10244 12782 10272 13874
rect 10704 13530 10732 14350
rect 11898 13628 12206 13648
rect 11898 13626 11904 13628
rect 11960 13626 11984 13628
rect 12040 13626 12064 13628
rect 12120 13626 12144 13628
rect 12200 13626 12206 13628
rect 11960 13574 11962 13626
rect 12142 13574 12144 13626
rect 11898 13572 11904 13574
rect 11960 13572 11984 13574
rect 12040 13572 12064 13574
rect 12120 13572 12144 13574
rect 12200 13572 12206 13574
rect 11898 13552 12206 13572
rect 10692 13524 10744 13530
rect 10692 13466 10744 13472
rect 10334 13084 10642 13104
rect 10334 13082 10340 13084
rect 10396 13082 10420 13084
rect 10476 13082 10500 13084
rect 10556 13082 10580 13084
rect 10636 13082 10642 13084
rect 10396 13030 10398 13082
rect 10578 13030 10580 13082
rect 10334 13028 10340 13030
rect 10396 13028 10420 13030
rect 10476 13028 10500 13030
rect 10556 13028 10580 13030
rect 10636 13028 10642 13030
rect 10334 13008 10642 13028
rect 10704 12986 10732 13466
rect 10968 13252 11020 13258
rect 10968 13194 11020 13200
rect 10692 12980 10744 12986
rect 10692 12922 10744 12928
rect 10140 12776 10192 12782
rect 10140 12718 10192 12724
rect 10232 12776 10284 12782
rect 10232 12718 10284 12724
rect 10048 12096 10100 12102
rect 10048 12038 10100 12044
rect 9680 11824 9732 11830
rect 9680 11766 9732 11772
rect 9588 11552 9640 11558
rect 9588 11494 9640 11500
rect 9600 11218 9628 11494
rect 9588 11212 9640 11218
rect 9588 11154 9640 11160
rect 9692 11150 9720 11766
rect 9680 11144 9732 11150
rect 9680 11086 9732 11092
rect 10152 10742 10180 12718
rect 10980 12714 11008 13194
rect 10968 12708 11020 12714
rect 10968 12650 11020 12656
rect 10980 12238 11008 12650
rect 11898 12540 12206 12560
rect 11898 12538 11904 12540
rect 11960 12538 11984 12540
rect 12040 12538 12064 12540
rect 12120 12538 12144 12540
rect 12200 12538 12206 12540
rect 11960 12486 11962 12538
rect 12142 12486 12144 12538
rect 11898 12484 11904 12486
rect 11960 12484 11984 12486
rect 12040 12484 12064 12486
rect 12120 12484 12144 12486
rect 12200 12484 12206 12486
rect 11898 12464 12206 12484
rect 10968 12232 11020 12238
rect 10968 12174 11020 12180
rect 10334 11996 10642 12016
rect 10334 11994 10340 11996
rect 10396 11994 10420 11996
rect 10476 11994 10500 11996
rect 10556 11994 10580 11996
rect 10636 11994 10642 11996
rect 10396 11942 10398 11994
rect 10578 11942 10580 11994
rect 10334 11940 10340 11942
rect 10396 11940 10420 11942
rect 10476 11940 10500 11942
rect 10556 11940 10580 11942
rect 10636 11940 10642 11942
rect 10334 11920 10642 11940
rect 10980 11830 11008 12174
rect 11336 12096 11388 12102
rect 11336 12038 11388 12044
rect 10968 11824 11020 11830
rect 10968 11766 11020 11772
rect 11348 11218 11376 12038
rect 11898 11452 12206 11472
rect 11898 11450 11904 11452
rect 11960 11450 11984 11452
rect 12040 11450 12064 11452
rect 12120 11450 12144 11452
rect 12200 11450 12206 11452
rect 11960 11398 11962 11450
rect 12142 11398 12144 11450
rect 11898 11396 11904 11398
rect 11960 11396 11984 11398
rect 12040 11396 12064 11398
rect 12120 11396 12144 11398
rect 12200 11396 12206 11398
rect 11898 11376 12206 11396
rect 11336 11212 11388 11218
rect 11336 11154 11388 11160
rect 10334 10908 10642 10928
rect 10334 10906 10340 10908
rect 10396 10906 10420 10908
rect 10476 10906 10500 10908
rect 10556 10906 10580 10908
rect 10636 10906 10642 10908
rect 10396 10854 10398 10906
rect 10578 10854 10580 10906
rect 10334 10852 10340 10854
rect 10396 10852 10420 10854
rect 10476 10852 10500 10854
rect 10556 10852 10580 10854
rect 10636 10852 10642 10854
rect 10334 10832 10642 10852
rect 10140 10736 10192 10742
rect 10140 10678 10192 10684
rect 9128 10668 9180 10674
rect 9128 10610 9180 10616
rect 9956 10668 10008 10674
rect 9956 10610 10008 10616
rect 10416 10668 10468 10674
rect 10416 10610 10468 10616
rect 8770 10364 9078 10384
rect 8770 10362 8776 10364
rect 8832 10362 8856 10364
rect 8912 10362 8936 10364
rect 8992 10362 9016 10364
rect 9072 10362 9078 10364
rect 8832 10310 8834 10362
rect 9014 10310 9016 10362
rect 8770 10308 8776 10310
rect 8832 10308 8856 10310
rect 8912 10308 8936 10310
rect 8992 10308 9016 10310
rect 9072 10308 9078 10310
rect 8770 10288 9078 10308
rect 9140 10146 9168 10610
rect 9772 10464 9824 10470
rect 9772 10406 9824 10412
rect 9048 10118 9168 10146
rect 9784 10130 9812 10406
rect 9772 10124 9824 10130
rect 9048 9518 9076 10118
rect 9772 10066 9824 10072
rect 9496 10056 9548 10062
rect 9496 9998 9548 10004
rect 9312 9580 9364 9586
rect 9312 9522 9364 9528
rect 9036 9512 9088 9518
rect 9036 9454 9088 9460
rect 8770 9276 9078 9296
rect 8770 9274 8776 9276
rect 8832 9274 8856 9276
rect 8912 9274 8936 9276
rect 8992 9274 9016 9276
rect 9072 9274 9078 9276
rect 8832 9222 8834 9274
rect 9014 9222 9016 9274
rect 8770 9220 8776 9222
rect 8832 9220 8856 9222
rect 8912 9220 8936 9222
rect 8992 9220 9016 9222
rect 9072 9220 9078 9222
rect 8770 9200 9078 9220
rect 9128 8492 9180 8498
rect 9128 8434 9180 8440
rect 8770 8188 9078 8208
rect 8770 8186 8776 8188
rect 8832 8186 8856 8188
rect 8912 8186 8936 8188
rect 8992 8186 9016 8188
rect 9072 8186 9078 8188
rect 8832 8134 8834 8186
rect 9014 8134 9016 8186
rect 8770 8132 8776 8134
rect 8832 8132 8856 8134
rect 8912 8132 8936 8134
rect 8992 8132 9016 8134
rect 9072 8132 9078 8134
rect 8770 8112 9078 8132
rect 9140 7970 9168 8434
rect 8956 7942 9168 7970
rect 8956 7886 8984 7942
rect 8300 7880 8352 7886
rect 8300 7822 8352 7828
rect 8944 7880 8996 7886
rect 8944 7822 8996 7828
rect 8300 7404 8352 7410
rect 8300 7346 8352 7352
rect 8312 6730 8340 7346
rect 8956 7342 8984 7822
rect 8944 7336 8996 7342
rect 8944 7278 8996 7284
rect 8770 7100 9078 7120
rect 8770 7098 8776 7100
rect 8832 7098 8856 7100
rect 8912 7098 8936 7100
rect 8992 7098 9016 7100
rect 9072 7098 9078 7100
rect 8832 7046 8834 7098
rect 9014 7046 9016 7098
rect 8770 7044 8776 7046
rect 8832 7044 8856 7046
rect 8912 7044 8936 7046
rect 8992 7044 9016 7046
rect 9072 7044 9078 7046
rect 8770 7024 9078 7044
rect 9324 6798 9352 9522
rect 9508 8974 9536 9998
rect 9968 9450 9996 10610
rect 10428 10130 10456 10610
rect 11898 10364 12206 10384
rect 11898 10362 11904 10364
rect 11960 10362 11984 10364
rect 12040 10362 12064 10364
rect 12120 10362 12144 10364
rect 12200 10362 12206 10364
rect 11960 10310 11962 10362
rect 12142 10310 12144 10362
rect 11898 10308 11904 10310
rect 11960 10308 11984 10310
rect 12040 10308 12064 10310
rect 12120 10308 12144 10310
rect 12200 10308 12206 10310
rect 11898 10288 12206 10308
rect 10416 10124 10468 10130
rect 10416 10066 10468 10072
rect 12452 10062 12480 14350
rect 12992 13320 13044 13326
rect 12992 13262 13044 13268
rect 12808 13184 12860 13190
rect 12808 13126 12860 13132
rect 12820 13025 12848 13126
rect 12806 13016 12862 13025
rect 12806 12951 12862 12960
rect 12716 12844 12768 12850
rect 12716 12786 12768 12792
rect 12728 11082 12756 12786
rect 12808 12776 12860 12782
rect 12808 12718 12860 12724
rect 12820 11354 12848 12718
rect 12808 11348 12860 11354
rect 12808 11290 12860 11296
rect 12716 11076 12768 11082
rect 12716 11018 12768 11024
rect 12624 10124 12676 10130
rect 12624 10066 12676 10072
rect 12440 10056 12492 10062
rect 12440 9998 12492 10004
rect 12164 9920 12216 9926
rect 12164 9862 12216 9868
rect 10334 9820 10642 9840
rect 10334 9818 10340 9820
rect 10396 9818 10420 9820
rect 10476 9818 10500 9820
rect 10556 9818 10580 9820
rect 10636 9818 10642 9820
rect 10396 9766 10398 9818
rect 10578 9766 10580 9818
rect 10334 9764 10340 9766
rect 10396 9764 10420 9766
rect 10476 9764 10500 9766
rect 10556 9764 10580 9766
rect 10636 9764 10642 9766
rect 10334 9744 10642 9764
rect 12176 9586 12204 9862
rect 12164 9580 12216 9586
rect 12164 9522 12216 9528
rect 9956 9444 10008 9450
rect 9956 9386 10008 9392
rect 11428 9376 11480 9382
rect 11428 9318 11480 9324
rect 11440 9042 11468 9318
rect 11898 9276 12206 9296
rect 11898 9274 11904 9276
rect 11960 9274 11984 9276
rect 12040 9274 12064 9276
rect 12120 9274 12144 9276
rect 12200 9274 12206 9276
rect 11960 9222 11962 9274
rect 12142 9222 12144 9274
rect 11898 9220 11904 9222
rect 11960 9220 11984 9222
rect 12040 9220 12064 9222
rect 12120 9220 12144 9222
rect 12200 9220 12206 9222
rect 11898 9200 12206 9220
rect 12452 9178 12480 9998
rect 12532 9920 12584 9926
rect 12532 9862 12584 9868
rect 12440 9172 12492 9178
rect 12440 9114 12492 9120
rect 11428 9036 11480 9042
rect 11428 8978 11480 8984
rect 9496 8968 9548 8974
rect 9496 8910 9548 8916
rect 10232 8968 10284 8974
rect 10232 8910 10284 8916
rect 9508 8634 9536 8910
rect 9496 8628 9548 8634
rect 9496 8570 9548 8576
rect 9496 7812 9548 7818
rect 9496 7754 9548 7760
rect 9508 7546 9536 7754
rect 9588 7744 9640 7750
rect 9588 7686 9640 7692
rect 9496 7540 9548 7546
rect 9496 7482 9548 7488
rect 9600 7478 9628 7686
rect 9588 7472 9640 7478
rect 9588 7414 9640 7420
rect 9600 7206 9628 7414
rect 9864 7336 9916 7342
rect 9864 7278 9916 7284
rect 9588 7200 9640 7206
rect 9588 7142 9640 7148
rect 9876 6934 9904 7278
rect 9864 6928 9916 6934
rect 9864 6870 9916 6876
rect 8576 6792 8628 6798
rect 8576 6734 8628 6740
rect 9312 6792 9364 6798
rect 9312 6734 9364 6740
rect 8300 6724 8352 6730
rect 8300 6666 8352 6672
rect 8312 6458 8340 6666
rect 8300 6452 8352 6458
rect 8300 6394 8352 6400
rect 8116 5364 8168 5370
rect 8116 5306 8168 5312
rect 7564 5296 7616 5302
rect 7564 5238 7616 5244
rect 7206 4380 7514 4400
rect 7206 4378 7212 4380
rect 7268 4378 7292 4380
rect 7348 4378 7372 4380
rect 7428 4378 7452 4380
rect 7508 4378 7514 4380
rect 7268 4326 7270 4378
rect 7450 4326 7452 4378
rect 7206 4324 7212 4326
rect 7268 4324 7292 4326
rect 7348 4324 7372 4326
rect 7428 4324 7452 4326
rect 7508 4324 7514 4326
rect 7206 4304 7514 4324
rect 7564 4208 7616 4214
rect 7564 4150 7616 4156
rect 7012 4140 7064 4146
rect 7012 4082 7064 4088
rect 6552 3936 6604 3942
rect 6552 3878 6604 3884
rect 5642 3836 5950 3856
rect 5642 3834 5648 3836
rect 5704 3834 5728 3836
rect 5784 3834 5808 3836
rect 5864 3834 5888 3836
rect 5944 3834 5950 3836
rect 5704 3782 5706 3834
rect 5886 3782 5888 3834
rect 5642 3780 5648 3782
rect 5704 3780 5728 3782
rect 5784 3780 5808 3782
rect 5864 3780 5888 3782
rect 5944 3780 5950 3782
rect 5642 3760 5950 3780
rect 5368 3590 5488 3618
rect 5368 3126 5396 3590
rect 5448 3528 5500 3534
rect 5448 3470 5500 3476
rect 5356 3120 5408 3126
rect 5356 3062 5408 3068
rect 4712 2984 4764 2990
rect 4712 2926 4764 2932
rect 5460 2650 5488 3470
rect 6368 3460 6420 3466
rect 6368 3402 6420 3408
rect 6380 3194 6408 3402
rect 6368 3188 6420 3194
rect 6368 3130 6420 3136
rect 6564 3058 6592 3878
rect 7576 3738 7604 4150
rect 8128 4146 8156 5306
rect 8588 4146 8616 6734
rect 8770 6012 9078 6032
rect 8770 6010 8776 6012
rect 8832 6010 8856 6012
rect 8912 6010 8936 6012
rect 8992 6010 9016 6012
rect 9072 6010 9078 6012
rect 8832 5958 8834 6010
rect 9014 5958 9016 6010
rect 8770 5956 8776 5958
rect 8832 5956 8856 5958
rect 8912 5956 8936 5958
rect 8992 5956 9016 5958
rect 9072 5956 9078 5958
rect 8770 5936 9078 5956
rect 9680 5772 9732 5778
rect 9680 5714 9732 5720
rect 9588 5364 9640 5370
rect 9588 5306 9640 5312
rect 9312 5296 9364 5302
rect 9312 5238 9364 5244
rect 8668 5160 8720 5166
rect 8668 5102 8720 5108
rect 9220 5160 9272 5166
rect 9220 5102 9272 5108
rect 8680 4690 8708 5102
rect 8770 4924 9078 4944
rect 8770 4922 8776 4924
rect 8832 4922 8856 4924
rect 8912 4922 8936 4924
rect 8992 4922 9016 4924
rect 9072 4922 9078 4924
rect 8832 4870 8834 4922
rect 9014 4870 9016 4922
rect 8770 4868 8776 4870
rect 8832 4868 8856 4870
rect 8912 4868 8936 4870
rect 8992 4868 9016 4870
rect 9072 4868 9078 4870
rect 8770 4848 9078 4868
rect 9232 4690 9260 5102
rect 8668 4684 8720 4690
rect 8668 4626 8720 4632
rect 9220 4684 9272 4690
rect 9220 4626 9272 4632
rect 8680 4214 8708 4626
rect 9324 4570 9352 5238
rect 9600 5234 9628 5306
rect 9692 5302 9720 5714
rect 9876 5710 9904 6870
rect 10244 6866 10272 8910
rect 10334 8732 10642 8752
rect 10334 8730 10340 8732
rect 10396 8730 10420 8732
rect 10476 8730 10500 8732
rect 10556 8730 10580 8732
rect 10636 8730 10642 8732
rect 10396 8678 10398 8730
rect 10578 8678 10580 8730
rect 10334 8676 10340 8678
rect 10396 8676 10420 8678
rect 10476 8676 10500 8678
rect 10556 8676 10580 8678
rect 10636 8676 10642 8678
rect 10334 8656 10642 8676
rect 11898 8188 12206 8208
rect 11898 8186 11904 8188
rect 11960 8186 11984 8188
rect 12040 8186 12064 8188
rect 12120 8186 12144 8188
rect 12200 8186 12206 8188
rect 11960 8134 11962 8186
rect 12142 8134 12144 8186
rect 11898 8132 11904 8134
rect 11960 8132 11984 8134
rect 12040 8132 12064 8134
rect 12120 8132 12144 8134
rect 12200 8132 12206 8134
rect 11898 8112 12206 8132
rect 12348 7812 12400 7818
rect 12348 7754 12400 7760
rect 10692 7744 10744 7750
rect 10692 7686 10744 7692
rect 10334 7644 10642 7664
rect 10334 7642 10340 7644
rect 10396 7642 10420 7644
rect 10476 7642 10500 7644
rect 10556 7642 10580 7644
rect 10636 7642 10642 7644
rect 10396 7590 10398 7642
rect 10578 7590 10580 7642
rect 10334 7588 10340 7590
rect 10396 7588 10420 7590
rect 10476 7588 10500 7590
rect 10556 7588 10580 7590
rect 10636 7588 10642 7590
rect 10334 7568 10642 7588
rect 10704 7342 10732 7686
rect 10968 7540 11020 7546
rect 10968 7482 11020 7488
rect 10692 7336 10744 7342
rect 10692 7278 10744 7284
rect 10980 6882 11008 7482
rect 11898 7100 12206 7120
rect 11898 7098 11904 7100
rect 11960 7098 11984 7100
rect 12040 7098 12064 7100
rect 12120 7098 12144 7100
rect 12200 7098 12206 7100
rect 11960 7046 11962 7098
rect 12142 7046 12144 7098
rect 11898 7044 11904 7046
rect 11960 7044 11984 7046
rect 12040 7044 12064 7046
rect 12120 7044 12144 7046
rect 12200 7044 12206 7046
rect 11898 7024 12206 7044
rect 10888 6866 11008 6882
rect 12360 6866 12388 7754
rect 10232 6860 10284 6866
rect 10232 6802 10284 6808
rect 10876 6860 11008 6866
rect 10928 6854 11008 6860
rect 12348 6860 12400 6866
rect 10876 6802 10928 6808
rect 12348 6802 12400 6808
rect 10334 6556 10642 6576
rect 10334 6554 10340 6556
rect 10396 6554 10420 6556
rect 10476 6554 10500 6556
rect 10556 6554 10580 6556
rect 10636 6554 10642 6556
rect 10396 6502 10398 6554
rect 10578 6502 10580 6554
rect 10334 6500 10340 6502
rect 10396 6500 10420 6502
rect 10476 6500 10500 6502
rect 10556 6500 10580 6502
rect 10636 6500 10642 6502
rect 10334 6480 10642 6500
rect 11898 6012 12206 6032
rect 11898 6010 11904 6012
rect 11960 6010 11984 6012
rect 12040 6010 12064 6012
rect 12120 6010 12144 6012
rect 12200 6010 12206 6012
rect 11960 5958 11962 6010
rect 12142 5958 12144 6010
rect 11898 5956 11904 5958
rect 11960 5956 11984 5958
rect 12040 5956 12064 5958
rect 12120 5956 12144 5958
rect 12200 5956 12206 5958
rect 11898 5936 12206 5956
rect 12544 5710 12572 9862
rect 12636 8498 12664 10066
rect 12728 9994 12756 11018
rect 12820 10130 12848 11290
rect 12808 10124 12860 10130
rect 12808 10066 12860 10072
rect 12716 9988 12768 9994
rect 12716 9930 12768 9936
rect 12728 8906 12756 9930
rect 12806 8936 12862 8945
rect 12716 8900 12768 8906
rect 12806 8871 12862 8880
rect 12716 8842 12768 8848
rect 12624 8492 12676 8498
rect 12624 8434 12676 8440
rect 12728 7546 12756 8842
rect 12820 8634 12848 8871
rect 12900 8832 12952 8838
rect 12900 8774 12952 8780
rect 12808 8628 12860 8634
rect 12808 8570 12860 8576
rect 12912 7954 12940 8774
rect 12900 7948 12952 7954
rect 12900 7890 12952 7896
rect 12808 7744 12860 7750
rect 12808 7686 12860 7692
rect 12716 7540 12768 7546
rect 12716 7482 12768 7488
rect 12820 7410 12848 7686
rect 12808 7404 12860 7410
rect 12808 7346 12860 7352
rect 12820 6730 12848 7346
rect 12808 6724 12860 6730
rect 12808 6666 12860 6672
rect 12820 5846 12848 6666
rect 13004 6254 13032 13262
rect 12992 6248 13044 6254
rect 12992 6190 13044 6196
rect 12808 5840 12860 5846
rect 12808 5782 12860 5788
rect 9864 5704 9916 5710
rect 9864 5646 9916 5652
rect 11336 5704 11388 5710
rect 11336 5646 11388 5652
rect 12532 5704 12584 5710
rect 12532 5646 12584 5652
rect 12808 5704 12860 5710
rect 12808 5646 12860 5652
rect 10334 5468 10642 5488
rect 10334 5466 10340 5468
rect 10396 5466 10420 5468
rect 10476 5466 10500 5468
rect 10556 5466 10580 5468
rect 10636 5466 10642 5468
rect 10396 5414 10398 5466
rect 10578 5414 10580 5466
rect 10334 5412 10340 5414
rect 10396 5412 10420 5414
rect 10476 5412 10500 5414
rect 10556 5412 10580 5414
rect 10636 5412 10642 5414
rect 10334 5392 10642 5412
rect 11348 5370 11376 5646
rect 12624 5636 12676 5642
rect 12624 5578 12676 5584
rect 11428 5568 11480 5574
rect 11428 5510 11480 5516
rect 11336 5364 11388 5370
rect 11336 5306 11388 5312
rect 9680 5296 9732 5302
rect 9680 5238 9732 5244
rect 9588 5228 9640 5234
rect 9588 5170 9640 5176
rect 10692 5228 10744 5234
rect 10692 5170 10744 5176
rect 10704 4622 10732 5170
rect 10784 5024 10836 5030
rect 10784 4966 10836 4972
rect 9232 4554 9352 4570
rect 10232 4616 10284 4622
rect 10232 4558 10284 4564
rect 10692 4616 10744 4622
rect 10692 4558 10744 4564
rect 9220 4548 9352 4554
rect 9272 4542 9352 4548
rect 9220 4490 9272 4496
rect 9232 4282 9260 4490
rect 9220 4276 9272 4282
rect 9220 4218 9272 4224
rect 10244 4214 10272 4558
rect 10692 4480 10744 4486
rect 10692 4422 10744 4428
rect 10334 4380 10642 4400
rect 10334 4378 10340 4380
rect 10396 4378 10420 4380
rect 10476 4378 10500 4380
rect 10556 4378 10580 4380
rect 10636 4378 10642 4380
rect 10396 4326 10398 4378
rect 10578 4326 10580 4378
rect 10334 4324 10340 4326
rect 10396 4324 10420 4326
rect 10476 4324 10500 4326
rect 10556 4324 10580 4326
rect 10636 4324 10642 4326
rect 10334 4304 10642 4324
rect 10704 4214 10732 4422
rect 8668 4208 8720 4214
rect 8668 4150 8720 4156
rect 10232 4208 10284 4214
rect 10232 4150 10284 4156
rect 10692 4208 10744 4214
rect 10692 4150 10744 4156
rect 8116 4140 8168 4146
rect 8116 4082 8168 4088
rect 8576 4140 8628 4146
rect 8576 4082 8628 4088
rect 8680 4026 8708 4150
rect 8588 3998 8708 4026
rect 10692 4072 10744 4078
rect 10692 4014 10744 4020
rect 8588 3738 8616 3998
rect 8668 3936 8720 3942
rect 8668 3878 8720 3884
rect 7564 3732 7616 3738
rect 7564 3674 7616 3680
rect 8576 3732 8628 3738
rect 8576 3674 8628 3680
rect 7104 3392 7156 3398
rect 7104 3334 7156 3340
rect 7116 3126 7144 3334
rect 7206 3292 7514 3312
rect 7206 3290 7212 3292
rect 7268 3290 7292 3292
rect 7348 3290 7372 3292
rect 7428 3290 7452 3292
rect 7508 3290 7514 3292
rect 7268 3238 7270 3290
rect 7450 3238 7452 3290
rect 7206 3236 7212 3238
rect 7268 3236 7292 3238
rect 7348 3236 7372 3238
rect 7428 3236 7452 3238
rect 7508 3236 7514 3238
rect 7206 3216 7514 3236
rect 7104 3120 7156 3126
rect 7104 3062 7156 3068
rect 6552 3052 6604 3058
rect 6552 2994 6604 3000
rect 5642 2748 5950 2768
rect 5642 2746 5648 2748
rect 5704 2746 5728 2748
rect 5784 2746 5808 2748
rect 5864 2746 5888 2748
rect 5944 2746 5950 2748
rect 5704 2694 5706 2746
rect 5886 2694 5888 2746
rect 5642 2692 5648 2694
rect 5704 2692 5728 2694
rect 5784 2692 5808 2694
rect 5864 2692 5888 2694
rect 5944 2692 5950 2694
rect 5642 2672 5950 2692
rect 5448 2644 5500 2650
rect 5448 2586 5500 2592
rect 4436 2576 4488 2582
rect 4436 2518 4488 2524
rect 3240 2508 3292 2514
rect 3240 2450 3292 2456
rect 7576 2446 7604 3674
rect 8680 3602 8708 3878
rect 8770 3836 9078 3856
rect 8770 3834 8776 3836
rect 8832 3834 8856 3836
rect 8912 3834 8936 3836
rect 8992 3834 9016 3836
rect 9072 3834 9078 3836
rect 8832 3782 8834 3834
rect 9014 3782 9016 3834
rect 8770 3780 8776 3782
rect 8832 3780 8856 3782
rect 8912 3780 8936 3782
rect 8992 3780 9016 3782
rect 9072 3780 9078 3782
rect 8770 3760 9078 3780
rect 10704 3738 10732 4014
rect 10692 3732 10744 3738
rect 10692 3674 10744 3680
rect 8668 3596 8720 3602
rect 8668 3538 8720 3544
rect 10334 3292 10642 3312
rect 10334 3290 10340 3292
rect 10396 3290 10420 3292
rect 10476 3290 10500 3292
rect 10556 3290 10580 3292
rect 10636 3290 10642 3292
rect 10396 3238 10398 3290
rect 10578 3238 10580 3290
rect 10334 3236 10340 3238
rect 10396 3236 10420 3238
rect 10476 3236 10500 3238
rect 10556 3236 10580 3238
rect 10636 3236 10642 3238
rect 10334 3216 10642 3236
rect 8770 2748 9078 2768
rect 8770 2746 8776 2748
rect 8832 2746 8856 2748
rect 8912 2746 8936 2748
rect 8992 2746 9016 2748
rect 9072 2746 9078 2748
rect 8832 2694 8834 2746
rect 9014 2694 9016 2746
rect 8770 2692 8776 2694
rect 8832 2692 8856 2694
rect 8912 2692 8936 2694
rect 8992 2692 9016 2694
rect 9072 2692 9078 2694
rect 8770 2672 9078 2692
rect 10704 2446 10732 3674
rect 10796 3466 10824 4966
rect 11440 4690 11468 5510
rect 12636 5234 12664 5578
rect 12624 5228 12676 5234
rect 12624 5170 12676 5176
rect 12716 5160 12768 5166
rect 12716 5102 12768 5108
rect 11898 4924 12206 4944
rect 11898 4922 11904 4924
rect 11960 4922 11984 4924
rect 12040 4922 12064 4924
rect 12120 4922 12144 4924
rect 12200 4922 12206 4924
rect 11960 4870 11962 4922
rect 12142 4870 12144 4922
rect 11898 4868 11904 4870
rect 11960 4868 11984 4870
rect 12040 4868 12064 4870
rect 12120 4868 12144 4870
rect 12200 4868 12206 4870
rect 11898 4848 12206 4868
rect 11428 4684 11480 4690
rect 11428 4626 11480 4632
rect 11152 4616 11204 4622
rect 11152 4558 11204 4564
rect 11164 4282 11192 4558
rect 12728 4554 12756 5102
rect 12716 4548 12768 4554
rect 12716 4490 12768 4496
rect 12728 4282 12756 4490
rect 12820 4486 12848 5646
rect 12898 4856 12954 4865
rect 12898 4791 12954 4800
rect 12808 4480 12860 4486
rect 12808 4422 12860 4428
rect 11152 4276 11204 4282
rect 11152 4218 11204 4224
rect 12716 4276 12768 4282
rect 12716 4218 12768 4224
rect 11898 3836 12206 3856
rect 11898 3834 11904 3836
rect 11960 3834 11984 3836
rect 12040 3834 12064 3836
rect 12120 3834 12144 3836
rect 12200 3834 12206 3836
rect 11960 3782 11962 3834
rect 12142 3782 12144 3834
rect 11898 3780 11904 3782
rect 11960 3780 11984 3782
rect 12040 3780 12064 3782
rect 12120 3780 12144 3782
rect 12200 3780 12206 3782
rect 11898 3760 12206 3780
rect 10784 3460 10836 3466
rect 10784 3402 10836 3408
rect 11898 2748 12206 2768
rect 11898 2746 11904 2748
rect 11960 2746 11984 2748
rect 12040 2746 12064 2748
rect 12120 2746 12144 2748
rect 12200 2746 12206 2748
rect 11960 2694 11962 2746
rect 12142 2694 12144 2746
rect 11898 2692 11904 2694
rect 11960 2692 11984 2694
rect 12040 2692 12064 2694
rect 12120 2692 12144 2694
rect 12200 2692 12206 2694
rect 11898 2672 12206 2692
rect 12820 2446 12848 4422
rect 12912 4146 12940 4791
rect 12900 4140 12952 4146
rect 12900 4082 12952 4088
rect 3884 2440 3936 2446
rect 3884 2382 3936 2388
rect 7564 2440 7616 2446
rect 7564 2382 7616 2388
rect 10692 2440 10744 2446
rect 10692 2382 10744 2388
rect 12808 2440 12860 2446
rect 12808 2382 12860 2388
rect 20 2372 72 2378
rect 20 2314 72 2320
rect 32 800 60 2314
rect 3896 800 3924 2382
rect 7748 2304 7800 2310
rect 7748 2246 7800 2252
rect 11612 2304 11664 2310
rect 11612 2246 11664 2252
rect 12348 2304 12400 2310
rect 12348 2246 12400 2252
rect 4078 2204 4386 2224
rect 4078 2202 4084 2204
rect 4140 2202 4164 2204
rect 4220 2202 4244 2204
rect 4300 2202 4324 2204
rect 4380 2202 4386 2204
rect 4140 2150 4142 2202
rect 4322 2150 4324 2202
rect 4078 2148 4084 2150
rect 4140 2148 4164 2150
rect 4220 2148 4244 2150
rect 4300 2148 4324 2150
rect 4380 2148 4386 2150
rect 4078 2128 4386 2148
rect 7206 2204 7514 2224
rect 7206 2202 7212 2204
rect 7268 2202 7292 2204
rect 7348 2202 7372 2204
rect 7428 2202 7452 2204
rect 7508 2202 7514 2204
rect 7268 2150 7270 2202
rect 7450 2150 7452 2202
rect 7206 2148 7212 2150
rect 7268 2148 7292 2150
rect 7348 2148 7372 2150
rect 7428 2148 7452 2150
rect 7508 2148 7514 2150
rect 7206 2128 7514 2148
rect 7760 800 7788 2246
rect 10334 2204 10642 2224
rect 10334 2202 10340 2204
rect 10396 2202 10420 2204
rect 10476 2202 10500 2204
rect 10556 2202 10580 2204
rect 10636 2202 10642 2204
rect 10396 2150 10398 2202
rect 10578 2150 10580 2202
rect 10334 2148 10340 2150
rect 10396 2148 10420 2150
rect 10476 2148 10500 2150
rect 10556 2148 10580 2150
rect 10636 2148 10642 2150
rect 10334 2128 10642 2148
rect 11624 800 11652 2246
rect 18 0 74 800
rect 3882 0 3938 800
rect 7746 0 7802 800
rect 11610 0 11666 800
rect 12360 785 12388 2246
rect 12346 776 12402 785
rect 12346 711 12402 720
<< via2 >>
rect 1490 15680 1546 15736
rect 2520 14714 2576 14716
rect 2600 14714 2656 14716
rect 2680 14714 2736 14716
rect 2760 14714 2816 14716
rect 2520 14662 2566 14714
rect 2566 14662 2576 14714
rect 2600 14662 2630 14714
rect 2630 14662 2642 14714
rect 2642 14662 2656 14714
rect 2680 14662 2694 14714
rect 2694 14662 2706 14714
rect 2706 14662 2736 14714
rect 2760 14662 2770 14714
rect 2770 14662 2816 14714
rect 2520 14660 2576 14662
rect 2600 14660 2656 14662
rect 2680 14660 2736 14662
rect 2760 14660 2816 14662
rect 5648 14714 5704 14716
rect 5728 14714 5784 14716
rect 5808 14714 5864 14716
rect 5888 14714 5944 14716
rect 5648 14662 5694 14714
rect 5694 14662 5704 14714
rect 5728 14662 5758 14714
rect 5758 14662 5770 14714
rect 5770 14662 5784 14714
rect 5808 14662 5822 14714
rect 5822 14662 5834 14714
rect 5834 14662 5864 14714
rect 5888 14662 5898 14714
rect 5898 14662 5944 14714
rect 5648 14660 5704 14662
rect 5728 14660 5784 14662
rect 5808 14660 5864 14662
rect 5888 14660 5944 14662
rect 8776 14714 8832 14716
rect 8856 14714 8912 14716
rect 8936 14714 8992 14716
rect 9016 14714 9072 14716
rect 8776 14662 8822 14714
rect 8822 14662 8832 14714
rect 8856 14662 8886 14714
rect 8886 14662 8898 14714
rect 8898 14662 8912 14714
rect 8936 14662 8950 14714
rect 8950 14662 8962 14714
rect 8962 14662 8992 14714
rect 9016 14662 9026 14714
rect 9026 14662 9072 14714
rect 8776 14660 8832 14662
rect 8856 14660 8912 14662
rect 8936 14660 8992 14662
rect 9016 14660 9072 14662
rect 11904 14714 11960 14716
rect 11984 14714 12040 14716
rect 12064 14714 12120 14716
rect 12144 14714 12200 14716
rect 11904 14662 11950 14714
rect 11950 14662 11960 14714
rect 11984 14662 12014 14714
rect 12014 14662 12026 14714
rect 12026 14662 12040 14714
rect 12064 14662 12078 14714
rect 12078 14662 12090 14714
rect 12090 14662 12120 14714
rect 12144 14662 12154 14714
rect 12154 14662 12200 14714
rect 11904 14660 11960 14662
rect 11984 14660 12040 14662
rect 12064 14660 12120 14662
rect 12144 14660 12200 14662
rect 2520 13626 2576 13628
rect 2600 13626 2656 13628
rect 2680 13626 2736 13628
rect 2760 13626 2816 13628
rect 2520 13574 2566 13626
rect 2566 13574 2576 13626
rect 2600 13574 2630 13626
rect 2630 13574 2642 13626
rect 2642 13574 2656 13626
rect 2680 13574 2694 13626
rect 2694 13574 2706 13626
rect 2706 13574 2736 13626
rect 2760 13574 2770 13626
rect 2770 13574 2816 13626
rect 2520 13572 2576 13574
rect 2600 13572 2656 13574
rect 2680 13572 2736 13574
rect 2760 13572 2816 13574
rect 2520 12538 2576 12540
rect 2600 12538 2656 12540
rect 2680 12538 2736 12540
rect 2760 12538 2816 12540
rect 2520 12486 2566 12538
rect 2566 12486 2576 12538
rect 2600 12486 2630 12538
rect 2630 12486 2642 12538
rect 2642 12486 2656 12538
rect 2680 12486 2694 12538
rect 2694 12486 2706 12538
rect 2706 12486 2736 12538
rect 2760 12486 2770 12538
rect 2770 12486 2816 12538
rect 2520 12484 2576 12486
rect 2600 12484 2656 12486
rect 2680 12484 2736 12486
rect 2760 12484 2816 12486
rect 1490 11620 1546 11656
rect 1490 11600 1492 11620
rect 1492 11600 1544 11620
rect 1544 11600 1546 11620
rect 1490 7520 1546 7576
rect 2520 11450 2576 11452
rect 2600 11450 2656 11452
rect 2680 11450 2736 11452
rect 2760 11450 2816 11452
rect 2520 11398 2566 11450
rect 2566 11398 2576 11450
rect 2600 11398 2630 11450
rect 2630 11398 2642 11450
rect 2642 11398 2656 11450
rect 2680 11398 2694 11450
rect 2694 11398 2706 11450
rect 2706 11398 2736 11450
rect 2760 11398 2770 11450
rect 2770 11398 2816 11450
rect 2520 11396 2576 11398
rect 2600 11396 2656 11398
rect 2680 11396 2736 11398
rect 2760 11396 2816 11398
rect 2520 10362 2576 10364
rect 2600 10362 2656 10364
rect 2680 10362 2736 10364
rect 2760 10362 2816 10364
rect 2520 10310 2566 10362
rect 2566 10310 2576 10362
rect 2600 10310 2630 10362
rect 2630 10310 2642 10362
rect 2642 10310 2656 10362
rect 2680 10310 2694 10362
rect 2694 10310 2706 10362
rect 2706 10310 2736 10362
rect 2760 10310 2770 10362
rect 2770 10310 2816 10362
rect 2520 10308 2576 10310
rect 2600 10308 2656 10310
rect 2680 10308 2736 10310
rect 2760 10308 2816 10310
rect 2520 9274 2576 9276
rect 2600 9274 2656 9276
rect 2680 9274 2736 9276
rect 2760 9274 2816 9276
rect 2520 9222 2566 9274
rect 2566 9222 2576 9274
rect 2600 9222 2630 9274
rect 2630 9222 2642 9274
rect 2642 9222 2656 9274
rect 2680 9222 2694 9274
rect 2694 9222 2706 9274
rect 2706 9222 2736 9274
rect 2760 9222 2770 9274
rect 2770 9222 2816 9274
rect 2520 9220 2576 9222
rect 2600 9220 2656 9222
rect 2680 9220 2736 9222
rect 2760 9220 2816 9222
rect 4084 14170 4140 14172
rect 4164 14170 4220 14172
rect 4244 14170 4300 14172
rect 4324 14170 4380 14172
rect 4084 14118 4130 14170
rect 4130 14118 4140 14170
rect 4164 14118 4194 14170
rect 4194 14118 4206 14170
rect 4206 14118 4220 14170
rect 4244 14118 4258 14170
rect 4258 14118 4270 14170
rect 4270 14118 4300 14170
rect 4324 14118 4334 14170
rect 4334 14118 4380 14170
rect 4084 14116 4140 14118
rect 4164 14116 4220 14118
rect 4244 14116 4300 14118
rect 4324 14116 4380 14118
rect 4084 13082 4140 13084
rect 4164 13082 4220 13084
rect 4244 13082 4300 13084
rect 4324 13082 4380 13084
rect 4084 13030 4130 13082
rect 4130 13030 4140 13082
rect 4164 13030 4194 13082
rect 4194 13030 4206 13082
rect 4206 13030 4220 13082
rect 4244 13030 4258 13082
rect 4258 13030 4270 13082
rect 4270 13030 4300 13082
rect 4324 13030 4334 13082
rect 4334 13030 4380 13082
rect 4084 13028 4140 13030
rect 4164 13028 4220 13030
rect 4244 13028 4300 13030
rect 4324 13028 4380 13030
rect 5648 13626 5704 13628
rect 5728 13626 5784 13628
rect 5808 13626 5864 13628
rect 5888 13626 5944 13628
rect 5648 13574 5694 13626
rect 5694 13574 5704 13626
rect 5728 13574 5758 13626
rect 5758 13574 5770 13626
rect 5770 13574 5784 13626
rect 5808 13574 5822 13626
rect 5822 13574 5834 13626
rect 5834 13574 5864 13626
rect 5888 13574 5898 13626
rect 5898 13574 5944 13626
rect 5648 13572 5704 13574
rect 5728 13572 5784 13574
rect 5808 13572 5864 13574
rect 5888 13572 5944 13574
rect 4084 11994 4140 11996
rect 4164 11994 4220 11996
rect 4244 11994 4300 11996
rect 4324 11994 4380 11996
rect 4084 11942 4130 11994
rect 4130 11942 4140 11994
rect 4164 11942 4194 11994
rect 4194 11942 4206 11994
rect 4206 11942 4220 11994
rect 4244 11942 4258 11994
rect 4258 11942 4270 11994
rect 4270 11942 4300 11994
rect 4324 11942 4334 11994
rect 4334 11942 4380 11994
rect 4084 11940 4140 11942
rect 4164 11940 4220 11942
rect 4244 11940 4300 11942
rect 4324 11940 4380 11942
rect 4084 10906 4140 10908
rect 4164 10906 4220 10908
rect 4244 10906 4300 10908
rect 4324 10906 4380 10908
rect 4084 10854 4130 10906
rect 4130 10854 4140 10906
rect 4164 10854 4194 10906
rect 4194 10854 4206 10906
rect 4206 10854 4220 10906
rect 4244 10854 4258 10906
rect 4258 10854 4270 10906
rect 4270 10854 4300 10906
rect 4324 10854 4334 10906
rect 4334 10854 4380 10906
rect 4084 10852 4140 10854
rect 4164 10852 4220 10854
rect 4244 10852 4300 10854
rect 4324 10852 4380 10854
rect 5648 12538 5704 12540
rect 5728 12538 5784 12540
rect 5808 12538 5864 12540
rect 5888 12538 5944 12540
rect 5648 12486 5694 12538
rect 5694 12486 5704 12538
rect 5728 12486 5758 12538
rect 5758 12486 5770 12538
rect 5770 12486 5784 12538
rect 5808 12486 5822 12538
rect 5822 12486 5834 12538
rect 5834 12486 5864 12538
rect 5888 12486 5898 12538
rect 5898 12486 5944 12538
rect 5648 12484 5704 12486
rect 5728 12484 5784 12486
rect 5808 12484 5864 12486
rect 5888 12484 5944 12486
rect 5648 11450 5704 11452
rect 5728 11450 5784 11452
rect 5808 11450 5864 11452
rect 5888 11450 5944 11452
rect 5648 11398 5694 11450
rect 5694 11398 5704 11450
rect 5728 11398 5758 11450
rect 5758 11398 5770 11450
rect 5770 11398 5784 11450
rect 5808 11398 5822 11450
rect 5822 11398 5834 11450
rect 5834 11398 5864 11450
rect 5888 11398 5898 11450
rect 5898 11398 5944 11450
rect 5648 11396 5704 11398
rect 5728 11396 5784 11398
rect 5808 11396 5864 11398
rect 5888 11396 5944 11398
rect 5648 10362 5704 10364
rect 5728 10362 5784 10364
rect 5808 10362 5864 10364
rect 5888 10362 5944 10364
rect 5648 10310 5694 10362
rect 5694 10310 5704 10362
rect 5728 10310 5758 10362
rect 5758 10310 5770 10362
rect 5770 10310 5784 10362
rect 5808 10310 5822 10362
rect 5822 10310 5834 10362
rect 5834 10310 5864 10362
rect 5888 10310 5898 10362
rect 5898 10310 5944 10362
rect 5648 10308 5704 10310
rect 5728 10308 5784 10310
rect 5808 10308 5864 10310
rect 5888 10308 5944 10310
rect 4084 9818 4140 9820
rect 4164 9818 4220 9820
rect 4244 9818 4300 9820
rect 4324 9818 4380 9820
rect 4084 9766 4130 9818
rect 4130 9766 4140 9818
rect 4164 9766 4194 9818
rect 4194 9766 4206 9818
rect 4206 9766 4220 9818
rect 4244 9766 4258 9818
rect 4258 9766 4270 9818
rect 4270 9766 4300 9818
rect 4324 9766 4334 9818
rect 4334 9766 4380 9818
rect 4084 9764 4140 9766
rect 4164 9764 4220 9766
rect 4244 9764 4300 9766
rect 4324 9764 4380 9766
rect 2520 8186 2576 8188
rect 2600 8186 2656 8188
rect 2680 8186 2736 8188
rect 2760 8186 2816 8188
rect 2520 8134 2566 8186
rect 2566 8134 2576 8186
rect 2600 8134 2630 8186
rect 2630 8134 2642 8186
rect 2642 8134 2656 8186
rect 2680 8134 2694 8186
rect 2694 8134 2706 8186
rect 2706 8134 2736 8186
rect 2760 8134 2770 8186
rect 2770 8134 2816 8186
rect 2520 8132 2576 8134
rect 2600 8132 2656 8134
rect 2680 8132 2736 8134
rect 2760 8132 2816 8134
rect 2520 7098 2576 7100
rect 2600 7098 2656 7100
rect 2680 7098 2736 7100
rect 2760 7098 2816 7100
rect 2520 7046 2566 7098
rect 2566 7046 2576 7098
rect 2600 7046 2630 7098
rect 2630 7046 2642 7098
rect 2642 7046 2656 7098
rect 2680 7046 2694 7098
rect 2694 7046 2706 7098
rect 2706 7046 2736 7098
rect 2760 7046 2770 7098
rect 2770 7046 2816 7098
rect 2520 7044 2576 7046
rect 2600 7044 2656 7046
rect 2680 7044 2736 7046
rect 2760 7044 2816 7046
rect 4084 8730 4140 8732
rect 4164 8730 4220 8732
rect 4244 8730 4300 8732
rect 4324 8730 4380 8732
rect 4084 8678 4130 8730
rect 4130 8678 4140 8730
rect 4164 8678 4194 8730
rect 4194 8678 4206 8730
rect 4206 8678 4220 8730
rect 4244 8678 4258 8730
rect 4258 8678 4270 8730
rect 4270 8678 4300 8730
rect 4324 8678 4334 8730
rect 4334 8678 4380 8730
rect 4084 8676 4140 8678
rect 4164 8676 4220 8678
rect 4244 8676 4300 8678
rect 4324 8676 4380 8678
rect 2520 6010 2576 6012
rect 2600 6010 2656 6012
rect 2680 6010 2736 6012
rect 2760 6010 2816 6012
rect 2520 5958 2566 6010
rect 2566 5958 2576 6010
rect 2600 5958 2630 6010
rect 2630 5958 2642 6010
rect 2642 5958 2656 6010
rect 2680 5958 2694 6010
rect 2694 5958 2706 6010
rect 2706 5958 2736 6010
rect 2760 5958 2770 6010
rect 2770 5958 2816 6010
rect 2520 5956 2576 5958
rect 2600 5956 2656 5958
rect 2680 5956 2736 5958
rect 2760 5956 2816 5958
rect 2520 4922 2576 4924
rect 2600 4922 2656 4924
rect 2680 4922 2736 4924
rect 2760 4922 2816 4924
rect 2520 4870 2566 4922
rect 2566 4870 2576 4922
rect 2600 4870 2630 4922
rect 2630 4870 2642 4922
rect 2642 4870 2656 4922
rect 2680 4870 2694 4922
rect 2694 4870 2706 4922
rect 2706 4870 2736 4922
rect 2760 4870 2770 4922
rect 2770 4870 2816 4922
rect 2520 4868 2576 4870
rect 2600 4868 2656 4870
rect 2680 4868 2736 4870
rect 2760 4868 2816 4870
rect 2520 3834 2576 3836
rect 2600 3834 2656 3836
rect 2680 3834 2736 3836
rect 2760 3834 2816 3836
rect 2520 3782 2566 3834
rect 2566 3782 2576 3834
rect 2600 3782 2630 3834
rect 2630 3782 2642 3834
rect 2642 3782 2656 3834
rect 2680 3782 2694 3834
rect 2694 3782 2706 3834
rect 2706 3782 2736 3834
rect 2760 3782 2770 3834
rect 2770 3782 2816 3834
rect 2520 3780 2576 3782
rect 2600 3780 2656 3782
rect 2680 3780 2736 3782
rect 2760 3780 2816 3782
rect 1490 3440 1546 3496
rect 2520 2746 2576 2748
rect 2600 2746 2656 2748
rect 2680 2746 2736 2748
rect 2760 2746 2816 2748
rect 2520 2694 2566 2746
rect 2566 2694 2576 2746
rect 2600 2694 2630 2746
rect 2630 2694 2642 2746
rect 2642 2694 2656 2746
rect 2680 2694 2694 2746
rect 2694 2694 2706 2746
rect 2706 2694 2736 2746
rect 2760 2694 2770 2746
rect 2770 2694 2816 2746
rect 2520 2692 2576 2694
rect 2600 2692 2656 2694
rect 2680 2692 2736 2694
rect 2760 2692 2816 2694
rect 4084 7642 4140 7644
rect 4164 7642 4220 7644
rect 4244 7642 4300 7644
rect 4324 7642 4380 7644
rect 4084 7590 4130 7642
rect 4130 7590 4140 7642
rect 4164 7590 4194 7642
rect 4194 7590 4206 7642
rect 4206 7590 4220 7642
rect 4244 7590 4258 7642
rect 4258 7590 4270 7642
rect 4270 7590 4300 7642
rect 4324 7590 4334 7642
rect 4334 7590 4380 7642
rect 4084 7588 4140 7590
rect 4164 7588 4220 7590
rect 4244 7588 4300 7590
rect 4324 7588 4380 7590
rect 4084 6554 4140 6556
rect 4164 6554 4220 6556
rect 4244 6554 4300 6556
rect 4324 6554 4380 6556
rect 4084 6502 4130 6554
rect 4130 6502 4140 6554
rect 4164 6502 4194 6554
rect 4194 6502 4206 6554
rect 4206 6502 4220 6554
rect 4244 6502 4258 6554
rect 4258 6502 4270 6554
rect 4270 6502 4300 6554
rect 4324 6502 4334 6554
rect 4334 6502 4380 6554
rect 4084 6500 4140 6502
rect 4164 6500 4220 6502
rect 4244 6500 4300 6502
rect 4324 6500 4380 6502
rect 5648 9274 5704 9276
rect 5728 9274 5784 9276
rect 5808 9274 5864 9276
rect 5888 9274 5944 9276
rect 5648 9222 5694 9274
rect 5694 9222 5704 9274
rect 5728 9222 5758 9274
rect 5758 9222 5770 9274
rect 5770 9222 5784 9274
rect 5808 9222 5822 9274
rect 5822 9222 5834 9274
rect 5834 9222 5864 9274
rect 5888 9222 5898 9274
rect 5898 9222 5944 9274
rect 5648 9220 5704 9222
rect 5728 9220 5784 9222
rect 5808 9220 5864 9222
rect 5888 9220 5944 9222
rect 5648 8186 5704 8188
rect 5728 8186 5784 8188
rect 5808 8186 5864 8188
rect 5888 8186 5944 8188
rect 5648 8134 5694 8186
rect 5694 8134 5704 8186
rect 5728 8134 5758 8186
rect 5758 8134 5770 8186
rect 5770 8134 5784 8186
rect 5808 8134 5822 8186
rect 5822 8134 5834 8186
rect 5834 8134 5864 8186
rect 5888 8134 5898 8186
rect 5898 8134 5944 8186
rect 5648 8132 5704 8134
rect 5728 8132 5784 8134
rect 5808 8132 5864 8134
rect 5888 8132 5944 8134
rect 7212 14170 7268 14172
rect 7292 14170 7348 14172
rect 7372 14170 7428 14172
rect 7452 14170 7508 14172
rect 7212 14118 7258 14170
rect 7258 14118 7268 14170
rect 7292 14118 7322 14170
rect 7322 14118 7334 14170
rect 7334 14118 7348 14170
rect 7372 14118 7386 14170
rect 7386 14118 7398 14170
rect 7398 14118 7428 14170
rect 7452 14118 7462 14170
rect 7462 14118 7508 14170
rect 7212 14116 7268 14118
rect 7292 14116 7348 14118
rect 7372 14116 7428 14118
rect 7452 14116 7508 14118
rect 10340 14170 10396 14172
rect 10420 14170 10476 14172
rect 10500 14170 10556 14172
rect 10580 14170 10636 14172
rect 10340 14118 10386 14170
rect 10386 14118 10396 14170
rect 10420 14118 10450 14170
rect 10450 14118 10462 14170
rect 10462 14118 10476 14170
rect 10500 14118 10514 14170
rect 10514 14118 10526 14170
rect 10526 14118 10556 14170
rect 10580 14118 10590 14170
rect 10590 14118 10636 14170
rect 10340 14116 10396 14118
rect 10420 14116 10476 14118
rect 10500 14116 10556 14118
rect 10580 14116 10636 14118
rect 8776 13626 8832 13628
rect 8856 13626 8912 13628
rect 8936 13626 8992 13628
rect 9016 13626 9072 13628
rect 8776 13574 8822 13626
rect 8822 13574 8832 13626
rect 8856 13574 8886 13626
rect 8886 13574 8898 13626
rect 8898 13574 8912 13626
rect 8936 13574 8950 13626
rect 8950 13574 8962 13626
rect 8962 13574 8992 13626
rect 9016 13574 9026 13626
rect 9026 13574 9072 13626
rect 8776 13572 8832 13574
rect 8856 13572 8912 13574
rect 8936 13572 8992 13574
rect 9016 13572 9072 13574
rect 7212 13082 7268 13084
rect 7292 13082 7348 13084
rect 7372 13082 7428 13084
rect 7452 13082 7508 13084
rect 7212 13030 7258 13082
rect 7258 13030 7268 13082
rect 7292 13030 7322 13082
rect 7322 13030 7334 13082
rect 7334 13030 7348 13082
rect 7372 13030 7386 13082
rect 7386 13030 7398 13082
rect 7398 13030 7428 13082
rect 7452 13030 7462 13082
rect 7462 13030 7508 13082
rect 7212 13028 7268 13030
rect 7292 13028 7348 13030
rect 7372 13028 7428 13030
rect 7452 13028 7508 13030
rect 7212 11994 7268 11996
rect 7292 11994 7348 11996
rect 7372 11994 7428 11996
rect 7452 11994 7508 11996
rect 7212 11942 7258 11994
rect 7258 11942 7268 11994
rect 7292 11942 7322 11994
rect 7322 11942 7334 11994
rect 7334 11942 7348 11994
rect 7372 11942 7386 11994
rect 7386 11942 7398 11994
rect 7398 11942 7428 11994
rect 7452 11942 7462 11994
rect 7462 11942 7508 11994
rect 7212 11940 7268 11942
rect 7292 11940 7348 11942
rect 7372 11940 7428 11942
rect 7452 11940 7508 11942
rect 7212 10906 7268 10908
rect 7292 10906 7348 10908
rect 7372 10906 7428 10908
rect 7452 10906 7508 10908
rect 7212 10854 7258 10906
rect 7258 10854 7268 10906
rect 7292 10854 7322 10906
rect 7322 10854 7334 10906
rect 7334 10854 7348 10906
rect 7372 10854 7386 10906
rect 7386 10854 7398 10906
rect 7398 10854 7428 10906
rect 7452 10854 7462 10906
rect 7462 10854 7508 10906
rect 7212 10852 7268 10854
rect 7292 10852 7348 10854
rect 7372 10852 7428 10854
rect 7452 10852 7508 10854
rect 8776 12538 8832 12540
rect 8856 12538 8912 12540
rect 8936 12538 8992 12540
rect 9016 12538 9072 12540
rect 8776 12486 8822 12538
rect 8822 12486 8832 12538
rect 8856 12486 8886 12538
rect 8886 12486 8898 12538
rect 8898 12486 8912 12538
rect 8936 12486 8950 12538
rect 8950 12486 8962 12538
rect 8962 12486 8992 12538
rect 9016 12486 9026 12538
rect 9026 12486 9072 12538
rect 8776 12484 8832 12486
rect 8856 12484 8912 12486
rect 8936 12484 8992 12486
rect 9016 12484 9072 12486
rect 8776 11450 8832 11452
rect 8856 11450 8912 11452
rect 8936 11450 8992 11452
rect 9016 11450 9072 11452
rect 8776 11398 8822 11450
rect 8822 11398 8832 11450
rect 8856 11398 8886 11450
rect 8886 11398 8898 11450
rect 8898 11398 8912 11450
rect 8936 11398 8950 11450
rect 8950 11398 8962 11450
rect 8962 11398 8992 11450
rect 9016 11398 9026 11450
rect 9026 11398 9072 11450
rect 8776 11396 8832 11398
rect 8856 11396 8912 11398
rect 8936 11396 8992 11398
rect 9016 11396 9072 11398
rect 7212 9818 7268 9820
rect 7292 9818 7348 9820
rect 7372 9818 7428 9820
rect 7452 9818 7508 9820
rect 7212 9766 7258 9818
rect 7258 9766 7268 9818
rect 7292 9766 7322 9818
rect 7322 9766 7334 9818
rect 7334 9766 7348 9818
rect 7372 9766 7386 9818
rect 7386 9766 7398 9818
rect 7398 9766 7428 9818
rect 7452 9766 7462 9818
rect 7462 9766 7508 9818
rect 7212 9764 7268 9766
rect 7292 9764 7348 9766
rect 7372 9764 7428 9766
rect 7452 9764 7508 9766
rect 7212 8730 7268 8732
rect 7292 8730 7348 8732
rect 7372 8730 7428 8732
rect 7452 8730 7508 8732
rect 7212 8678 7258 8730
rect 7258 8678 7268 8730
rect 7292 8678 7322 8730
rect 7322 8678 7334 8730
rect 7334 8678 7348 8730
rect 7372 8678 7386 8730
rect 7386 8678 7398 8730
rect 7398 8678 7428 8730
rect 7452 8678 7462 8730
rect 7462 8678 7508 8730
rect 7212 8676 7268 8678
rect 7292 8676 7348 8678
rect 7372 8676 7428 8678
rect 7452 8676 7508 8678
rect 5648 7098 5704 7100
rect 5728 7098 5784 7100
rect 5808 7098 5864 7100
rect 5888 7098 5944 7100
rect 5648 7046 5694 7098
rect 5694 7046 5704 7098
rect 5728 7046 5758 7098
rect 5758 7046 5770 7098
rect 5770 7046 5784 7098
rect 5808 7046 5822 7098
rect 5822 7046 5834 7098
rect 5834 7046 5864 7098
rect 5888 7046 5898 7098
rect 5898 7046 5944 7098
rect 5648 7044 5704 7046
rect 5728 7044 5784 7046
rect 5808 7044 5864 7046
rect 5888 7044 5944 7046
rect 7212 7642 7268 7644
rect 7292 7642 7348 7644
rect 7372 7642 7428 7644
rect 7452 7642 7508 7644
rect 7212 7590 7258 7642
rect 7258 7590 7268 7642
rect 7292 7590 7322 7642
rect 7322 7590 7334 7642
rect 7334 7590 7348 7642
rect 7372 7590 7386 7642
rect 7386 7590 7398 7642
rect 7398 7590 7428 7642
rect 7452 7590 7462 7642
rect 7462 7590 7508 7642
rect 7212 7588 7268 7590
rect 7292 7588 7348 7590
rect 7372 7588 7428 7590
rect 7452 7588 7508 7590
rect 4084 5466 4140 5468
rect 4164 5466 4220 5468
rect 4244 5466 4300 5468
rect 4324 5466 4380 5468
rect 4084 5414 4130 5466
rect 4130 5414 4140 5466
rect 4164 5414 4194 5466
rect 4194 5414 4206 5466
rect 4206 5414 4220 5466
rect 4244 5414 4258 5466
rect 4258 5414 4270 5466
rect 4270 5414 4300 5466
rect 4324 5414 4334 5466
rect 4334 5414 4380 5466
rect 4084 5412 4140 5414
rect 4164 5412 4220 5414
rect 4244 5412 4300 5414
rect 4324 5412 4380 5414
rect 4084 4378 4140 4380
rect 4164 4378 4220 4380
rect 4244 4378 4300 4380
rect 4324 4378 4380 4380
rect 4084 4326 4130 4378
rect 4130 4326 4140 4378
rect 4164 4326 4194 4378
rect 4194 4326 4206 4378
rect 4206 4326 4220 4378
rect 4244 4326 4258 4378
rect 4258 4326 4270 4378
rect 4270 4326 4300 4378
rect 4324 4326 4334 4378
rect 4334 4326 4380 4378
rect 4084 4324 4140 4326
rect 4164 4324 4220 4326
rect 4244 4324 4300 4326
rect 4324 4324 4380 4326
rect 4084 3290 4140 3292
rect 4164 3290 4220 3292
rect 4244 3290 4300 3292
rect 4324 3290 4380 3292
rect 4084 3238 4130 3290
rect 4130 3238 4140 3290
rect 4164 3238 4194 3290
rect 4194 3238 4206 3290
rect 4206 3238 4220 3290
rect 4244 3238 4258 3290
rect 4258 3238 4270 3290
rect 4270 3238 4300 3290
rect 4324 3238 4334 3290
rect 4334 3238 4380 3290
rect 4084 3236 4140 3238
rect 4164 3236 4220 3238
rect 4244 3236 4300 3238
rect 4324 3236 4380 3238
rect 5648 6010 5704 6012
rect 5728 6010 5784 6012
rect 5808 6010 5864 6012
rect 5888 6010 5944 6012
rect 5648 5958 5694 6010
rect 5694 5958 5704 6010
rect 5728 5958 5758 6010
rect 5758 5958 5770 6010
rect 5770 5958 5784 6010
rect 5808 5958 5822 6010
rect 5822 5958 5834 6010
rect 5834 5958 5864 6010
rect 5888 5958 5898 6010
rect 5898 5958 5944 6010
rect 5648 5956 5704 5958
rect 5728 5956 5784 5958
rect 5808 5956 5864 5958
rect 5888 5956 5944 5958
rect 5648 4922 5704 4924
rect 5728 4922 5784 4924
rect 5808 4922 5864 4924
rect 5888 4922 5944 4924
rect 5648 4870 5694 4922
rect 5694 4870 5704 4922
rect 5728 4870 5758 4922
rect 5758 4870 5770 4922
rect 5770 4870 5784 4922
rect 5808 4870 5822 4922
rect 5822 4870 5834 4922
rect 5834 4870 5864 4922
rect 5888 4870 5898 4922
rect 5898 4870 5944 4922
rect 5648 4868 5704 4870
rect 5728 4868 5784 4870
rect 5808 4868 5864 4870
rect 5888 4868 5944 4870
rect 7212 6554 7268 6556
rect 7292 6554 7348 6556
rect 7372 6554 7428 6556
rect 7452 6554 7508 6556
rect 7212 6502 7258 6554
rect 7258 6502 7268 6554
rect 7292 6502 7322 6554
rect 7322 6502 7334 6554
rect 7334 6502 7348 6554
rect 7372 6502 7386 6554
rect 7386 6502 7398 6554
rect 7398 6502 7428 6554
rect 7452 6502 7462 6554
rect 7462 6502 7508 6554
rect 7212 6500 7268 6502
rect 7292 6500 7348 6502
rect 7372 6500 7428 6502
rect 7452 6500 7508 6502
rect 7212 5466 7268 5468
rect 7292 5466 7348 5468
rect 7372 5466 7428 5468
rect 7452 5466 7508 5468
rect 7212 5414 7258 5466
rect 7258 5414 7268 5466
rect 7292 5414 7322 5466
rect 7322 5414 7334 5466
rect 7334 5414 7348 5466
rect 7372 5414 7386 5466
rect 7386 5414 7398 5466
rect 7398 5414 7428 5466
rect 7452 5414 7462 5466
rect 7462 5414 7508 5466
rect 7212 5412 7268 5414
rect 7292 5412 7348 5414
rect 7372 5412 7428 5414
rect 7452 5412 7508 5414
rect 11904 13626 11960 13628
rect 11984 13626 12040 13628
rect 12064 13626 12120 13628
rect 12144 13626 12200 13628
rect 11904 13574 11950 13626
rect 11950 13574 11960 13626
rect 11984 13574 12014 13626
rect 12014 13574 12026 13626
rect 12026 13574 12040 13626
rect 12064 13574 12078 13626
rect 12078 13574 12090 13626
rect 12090 13574 12120 13626
rect 12144 13574 12154 13626
rect 12154 13574 12200 13626
rect 11904 13572 11960 13574
rect 11984 13572 12040 13574
rect 12064 13572 12120 13574
rect 12144 13572 12200 13574
rect 10340 13082 10396 13084
rect 10420 13082 10476 13084
rect 10500 13082 10556 13084
rect 10580 13082 10636 13084
rect 10340 13030 10386 13082
rect 10386 13030 10396 13082
rect 10420 13030 10450 13082
rect 10450 13030 10462 13082
rect 10462 13030 10476 13082
rect 10500 13030 10514 13082
rect 10514 13030 10526 13082
rect 10526 13030 10556 13082
rect 10580 13030 10590 13082
rect 10590 13030 10636 13082
rect 10340 13028 10396 13030
rect 10420 13028 10476 13030
rect 10500 13028 10556 13030
rect 10580 13028 10636 13030
rect 11904 12538 11960 12540
rect 11984 12538 12040 12540
rect 12064 12538 12120 12540
rect 12144 12538 12200 12540
rect 11904 12486 11950 12538
rect 11950 12486 11960 12538
rect 11984 12486 12014 12538
rect 12014 12486 12026 12538
rect 12026 12486 12040 12538
rect 12064 12486 12078 12538
rect 12078 12486 12090 12538
rect 12090 12486 12120 12538
rect 12144 12486 12154 12538
rect 12154 12486 12200 12538
rect 11904 12484 11960 12486
rect 11984 12484 12040 12486
rect 12064 12484 12120 12486
rect 12144 12484 12200 12486
rect 10340 11994 10396 11996
rect 10420 11994 10476 11996
rect 10500 11994 10556 11996
rect 10580 11994 10636 11996
rect 10340 11942 10386 11994
rect 10386 11942 10396 11994
rect 10420 11942 10450 11994
rect 10450 11942 10462 11994
rect 10462 11942 10476 11994
rect 10500 11942 10514 11994
rect 10514 11942 10526 11994
rect 10526 11942 10556 11994
rect 10580 11942 10590 11994
rect 10590 11942 10636 11994
rect 10340 11940 10396 11942
rect 10420 11940 10476 11942
rect 10500 11940 10556 11942
rect 10580 11940 10636 11942
rect 11904 11450 11960 11452
rect 11984 11450 12040 11452
rect 12064 11450 12120 11452
rect 12144 11450 12200 11452
rect 11904 11398 11950 11450
rect 11950 11398 11960 11450
rect 11984 11398 12014 11450
rect 12014 11398 12026 11450
rect 12026 11398 12040 11450
rect 12064 11398 12078 11450
rect 12078 11398 12090 11450
rect 12090 11398 12120 11450
rect 12144 11398 12154 11450
rect 12154 11398 12200 11450
rect 11904 11396 11960 11398
rect 11984 11396 12040 11398
rect 12064 11396 12120 11398
rect 12144 11396 12200 11398
rect 10340 10906 10396 10908
rect 10420 10906 10476 10908
rect 10500 10906 10556 10908
rect 10580 10906 10636 10908
rect 10340 10854 10386 10906
rect 10386 10854 10396 10906
rect 10420 10854 10450 10906
rect 10450 10854 10462 10906
rect 10462 10854 10476 10906
rect 10500 10854 10514 10906
rect 10514 10854 10526 10906
rect 10526 10854 10556 10906
rect 10580 10854 10590 10906
rect 10590 10854 10636 10906
rect 10340 10852 10396 10854
rect 10420 10852 10476 10854
rect 10500 10852 10556 10854
rect 10580 10852 10636 10854
rect 8776 10362 8832 10364
rect 8856 10362 8912 10364
rect 8936 10362 8992 10364
rect 9016 10362 9072 10364
rect 8776 10310 8822 10362
rect 8822 10310 8832 10362
rect 8856 10310 8886 10362
rect 8886 10310 8898 10362
rect 8898 10310 8912 10362
rect 8936 10310 8950 10362
rect 8950 10310 8962 10362
rect 8962 10310 8992 10362
rect 9016 10310 9026 10362
rect 9026 10310 9072 10362
rect 8776 10308 8832 10310
rect 8856 10308 8912 10310
rect 8936 10308 8992 10310
rect 9016 10308 9072 10310
rect 8776 9274 8832 9276
rect 8856 9274 8912 9276
rect 8936 9274 8992 9276
rect 9016 9274 9072 9276
rect 8776 9222 8822 9274
rect 8822 9222 8832 9274
rect 8856 9222 8886 9274
rect 8886 9222 8898 9274
rect 8898 9222 8912 9274
rect 8936 9222 8950 9274
rect 8950 9222 8962 9274
rect 8962 9222 8992 9274
rect 9016 9222 9026 9274
rect 9026 9222 9072 9274
rect 8776 9220 8832 9222
rect 8856 9220 8912 9222
rect 8936 9220 8992 9222
rect 9016 9220 9072 9222
rect 8776 8186 8832 8188
rect 8856 8186 8912 8188
rect 8936 8186 8992 8188
rect 9016 8186 9072 8188
rect 8776 8134 8822 8186
rect 8822 8134 8832 8186
rect 8856 8134 8886 8186
rect 8886 8134 8898 8186
rect 8898 8134 8912 8186
rect 8936 8134 8950 8186
rect 8950 8134 8962 8186
rect 8962 8134 8992 8186
rect 9016 8134 9026 8186
rect 9026 8134 9072 8186
rect 8776 8132 8832 8134
rect 8856 8132 8912 8134
rect 8936 8132 8992 8134
rect 9016 8132 9072 8134
rect 8776 7098 8832 7100
rect 8856 7098 8912 7100
rect 8936 7098 8992 7100
rect 9016 7098 9072 7100
rect 8776 7046 8822 7098
rect 8822 7046 8832 7098
rect 8856 7046 8886 7098
rect 8886 7046 8898 7098
rect 8898 7046 8912 7098
rect 8936 7046 8950 7098
rect 8950 7046 8962 7098
rect 8962 7046 8992 7098
rect 9016 7046 9026 7098
rect 9026 7046 9072 7098
rect 8776 7044 8832 7046
rect 8856 7044 8912 7046
rect 8936 7044 8992 7046
rect 9016 7044 9072 7046
rect 11904 10362 11960 10364
rect 11984 10362 12040 10364
rect 12064 10362 12120 10364
rect 12144 10362 12200 10364
rect 11904 10310 11950 10362
rect 11950 10310 11960 10362
rect 11984 10310 12014 10362
rect 12014 10310 12026 10362
rect 12026 10310 12040 10362
rect 12064 10310 12078 10362
rect 12078 10310 12090 10362
rect 12090 10310 12120 10362
rect 12144 10310 12154 10362
rect 12154 10310 12200 10362
rect 11904 10308 11960 10310
rect 11984 10308 12040 10310
rect 12064 10308 12120 10310
rect 12144 10308 12200 10310
rect 12806 12960 12862 13016
rect 10340 9818 10396 9820
rect 10420 9818 10476 9820
rect 10500 9818 10556 9820
rect 10580 9818 10636 9820
rect 10340 9766 10386 9818
rect 10386 9766 10396 9818
rect 10420 9766 10450 9818
rect 10450 9766 10462 9818
rect 10462 9766 10476 9818
rect 10500 9766 10514 9818
rect 10514 9766 10526 9818
rect 10526 9766 10556 9818
rect 10580 9766 10590 9818
rect 10590 9766 10636 9818
rect 10340 9764 10396 9766
rect 10420 9764 10476 9766
rect 10500 9764 10556 9766
rect 10580 9764 10636 9766
rect 11904 9274 11960 9276
rect 11984 9274 12040 9276
rect 12064 9274 12120 9276
rect 12144 9274 12200 9276
rect 11904 9222 11950 9274
rect 11950 9222 11960 9274
rect 11984 9222 12014 9274
rect 12014 9222 12026 9274
rect 12026 9222 12040 9274
rect 12064 9222 12078 9274
rect 12078 9222 12090 9274
rect 12090 9222 12120 9274
rect 12144 9222 12154 9274
rect 12154 9222 12200 9274
rect 11904 9220 11960 9222
rect 11984 9220 12040 9222
rect 12064 9220 12120 9222
rect 12144 9220 12200 9222
rect 7212 4378 7268 4380
rect 7292 4378 7348 4380
rect 7372 4378 7428 4380
rect 7452 4378 7508 4380
rect 7212 4326 7258 4378
rect 7258 4326 7268 4378
rect 7292 4326 7322 4378
rect 7322 4326 7334 4378
rect 7334 4326 7348 4378
rect 7372 4326 7386 4378
rect 7386 4326 7398 4378
rect 7398 4326 7428 4378
rect 7452 4326 7462 4378
rect 7462 4326 7508 4378
rect 7212 4324 7268 4326
rect 7292 4324 7348 4326
rect 7372 4324 7428 4326
rect 7452 4324 7508 4326
rect 5648 3834 5704 3836
rect 5728 3834 5784 3836
rect 5808 3834 5864 3836
rect 5888 3834 5944 3836
rect 5648 3782 5694 3834
rect 5694 3782 5704 3834
rect 5728 3782 5758 3834
rect 5758 3782 5770 3834
rect 5770 3782 5784 3834
rect 5808 3782 5822 3834
rect 5822 3782 5834 3834
rect 5834 3782 5864 3834
rect 5888 3782 5898 3834
rect 5898 3782 5944 3834
rect 5648 3780 5704 3782
rect 5728 3780 5784 3782
rect 5808 3780 5864 3782
rect 5888 3780 5944 3782
rect 8776 6010 8832 6012
rect 8856 6010 8912 6012
rect 8936 6010 8992 6012
rect 9016 6010 9072 6012
rect 8776 5958 8822 6010
rect 8822 5958 8832 6010
rect 8856 5958 8886 6010
rect 8886 5958 8898 6010
rect 8898 5958 8912 6010
rect 8936 5958 8950 6010
rect 8950 5958 8962 6010
rect 8962 5958 8992 6010
rect 9016 5958 9026 6010
rect 9026 5958 9072 6010
rect 8776 5956 8832 5958
rect 8856 5956 8912 5958
rect 8936 5956 8992 5958
rect 9016 5956 9072 5958
rect 8776 4922 8832 4924
rect 8856 4922 8912 4924
rect 8936 4922 8992 4924
rect 9016 4922 9072 4924
rect 8776 4870 8822 4922
rect 8822 4870 8832 4922
rect 8856 4870 8886 4922
rect 8886 4870 8898 4922
rect 8898 4870 8912 4922
rect 8936 4870 8950 4922
rect 8950 4870 8962 4922
rect 8962 4870 8992 4922
rect 9016 4870 9026 4922
rect 9026 4870 9072 4922
rect 8776 4868 8832 4870
rect 8856 4868 8912 4870
rect 8936 4868 8992 4870
rect 9016 4868 9072 4870
rect 10340 8730 10396 8732
rect 10420 8730 10476 8732
rect 10500 8730 10556 8732
rect 10580 8730 10636 8732
rect 10340 8678 10386 8730
rect 10386 8678 10396 8730
rect 10420 8678 10450 8730
rect 10450 8678 10462 8730
rect 10462 8678 10476 8730
rect 10500 8678 10514 8730
rect 10514 8678 10526 8730
rect 10526 8678 10556 8730
rect 10580 8678 10590 8730
rect 10590 8678 10636 8730
rect 10340 8676 10396 8678
rect 10420 8676 10476 8678
rect 10500 8676 10556 8678
rect 10580 8676 10636 8678
rect 11904 8186 11960 8188
rect 11984 8186 12040 8188
rect 12064 8186 12120 8188
rect 12144 8186 12200 8188
rect 11904 8134 11950 8186
rect 11950 8134 11960 8186
rect 11984 8134 12014 8186
rect 12014 8134 12026 8186
rect 12026 8134 12040 8186
rect 12064 8134 12078 8186
rect 12078 8134 12090 8186
rect 12090 8134 12120 8186
rect 12144 8134 12154 8186
rect 12154 8134 12200 8186
rect 11904 8132 11960 8134
rect 11984 8132 12040 8134
rect 12064 8132 12120 8134
rect 12144 8132 12200 8134
rect 10340 7642 10396 7644
rect 10420 7642 10476 7644
rect 10500 7642 10556 7644
rect 10580 7642 10636 7644
rect 10340 7590 10386 7642
rect 10386 7590 10396 7642
rect 10420 7590 10450 7642
rect 10450 7590 10462 7642
rect 10462 7590 10476 7642
rect 10500 7590 10514 7642
rect 10514 7590 10526 7642
rect 10526 7590 10556 7642
rect 10580 7590 10590 7642
rect 10590 7590 10636 7642
rect 10340 7588 10396 7590
rect 10420 7588 10476 7590
rect 10500 7588 10556 7590
rect 10580 7588 10636 7590
rect 11904 7098 11960 7100
rect 11984 7098 12040 7100
rect 12064 7098 12120 7100
rect 12144 7098 12200 7100
rect 11904 7046 11950 7098
rect 11950 7046 11960 7098
rect 11984 7046 12014 7098
rect 12014 7046 12026 7098
rect 12026 7046 12040 7098
rect 12064 7046 12078 7098
rect 12078 7046 12090 7098
rect 12090 7046 12120 7098
rect 12144 7046 12154 7098
rect 12154 7046 12200 7098
rect 11904 7044 11960 7046
rect 11984 7044 12040 7046
rect 12064 7044 12120 7046
rect 12144 7044 12200 7046
rect 10340 6554 10396 6556
rect 10420 6554 10476 6556
rect 10500 6554 10556 6556
rect 10580 6554 10636 6556
rect 10340 6502 10386 6554
rect 10386 6502 10396 6554
rect 10420 6502 10450 6554
rect 10450 6502 10462 6554
rect 10462 6502 10476 6554
rect 10500 6502 10514 6554
rect 10514 6502 10526 6554
rect 10526 6502 10556 6554
rect 10580 6502 10590 6554
rect 10590 6502 10636 6554
rect 10340 6500 10396 6502
rect 10420 6500 10476 6502
rect 10500 6500 10556 6502
rect 10580 6500 10636 6502
rect 11904 6010 11960 6012
rect 11984 6010 12040 6012
rect 12064 6010 12120 6012
rect 12144 6010 12200 6012
rect 11904 5958 11950 6010
rect 11950 5958 11960 6010
rect 11984 5958 12014 6010
rect 12014 5958 12026 6010
rect 12026 5958 12040 6010
rect 12064 5958 12078 6010
rect 12078 5958 12090 6010
rect 12090 5958 12120 6010
rect 12144 5958 12154 6010
rect 12154 5958 12200 6010
rect 11904 5956 11960 5958
rect 11984 5956 12040 5958
rect 12064 5956 12120 5958
rect 12144 5956 12200 5958
rect 12806 8880 12862 8936
rect 10340 5466 10396 5468
rect 10420 5466 10476 5468
rect 10500 5466 10556 5468
rect 10580 5466 10636 5468
rect 10340 5414 10386 5466
rect 10386 5414 10396 5466
rect 10420 5414 10450 5466
rect 10450 5414 10462 5466
rect 10462 5414 10476 5466
rect 10500 5414 10514 5466
rect 10514 5414 10526 5466
rect 10526 5414 10556 5466
rect 10580 5414 10590 5466
rect 10590 5414 10636 5466
rect 10340 5412 10396 5414
rect 10420 5412 10476 5414
rect 10500 5412 10556 5414
rect 10580 5412 10636 5414
rect 10340 4378 10396 4380
rect 10420 4378 10476 4380
rect 10500 4378 10556 4380
rect 10580 4378 10636 4380
rect 10340 4326 10386 4378
rect 10386 4326 10396 4378
rect 10420 4326 10450 4378
rect 10450 4326 10462 4378
rect 10462 4326 10476 4378
rect 10500 4326 10514 4378
rect 10514 4326 10526 4378
rect 10526 4326 10556 4378
rect 10580 4326 10590 4378
rect 10590 4326 10636 4378
rect 10340 4324 10396 4326
rect 10420 4324 10476 4326
rect 10500 4324 10556 4326
rect 10580 4324 10636 4326
rect 7212 3290 7268 3292
rect 7292 3290 7348 3292
rect 7372 3290 7428 3292
rect 7452 3290 7508 3292
rect 7212 3238 7258 3290
rect 7258 3238 7268 3290
rect 7292 3238 7322 3290
rect 7322 3238 7334 3290
rect 7334 3238 7348 3290
rect 7372 3238 7386 3290
rect 7386 3238 7398 3290
rect 7398 3238 7428 3290
rect 7452 3238 7462 3290
rect 7462 3238 7508 3290
rect 7212 3236 7268 3238
rect 7292 3236 7348 3238
rect 7372 3236 7428 3238
rect 7452 3236 7508 3238
rect 5648 2746 5704 2748
rect 5728 2746 5784 2748
rect 5808 2746 5864 2748
rect 5888 2746 5944 2748
rect 5648 2694 5694 2746
rect 5694 2694 5704 2746
rect 5728 2694 5758 2746
rect 5758 2694 5770 2746
rect 5770 2694 5784 2746
rect 5808 2694 5822 2746
rect 5822 2694 5834 2746
rect 5834 2694 5864 2746
rect 5888 2694 5898 2746
rect 5898 2694 5944 2746
rect 5648 2692 5704 2694
rect 5728 2692 5784 2694
rect 5808 2692 5864 2694
rect 5888 2692 5944 2694
rect 8776 3834 8832 3836
rect 8856 3834 8912 3836
rect 8936 3834 8992 3836
rect 9016 3834 9072 3836
rect 8776 3782 8822 3834
rect 8822 3782 8832 3834
rect 8856 3782 8886 3834
rect 8886 3782 8898 3834
rect 8898 3782 8912 3834
rect 8936 3782 8950 3834
rect 8950 3782 8962 3834
rect 8962 3782 8992 3834
rect 9016 3782 9026 3834
rect 9026 3782 9072 3834
rect 8776 3780 8832 3782
rect 8856 3780 8912 3782
rect 8936 3780 8992 3782
rect 9016 3780 9072 3782
rect 10340 3290 10396 3292
rect 10420 3290 10476 3292
rect 10500 3290 10556 3292
rect 10580 3290 10636 3292
rect 10340 3238 10386 3290
rect 10386 3238 10396 3290
rect 10420 3238 10450 3290
rect 10450 3238 10462 3290
rect 10462 3238 10476 3290
rect 10500 3238 10514 3290
rect 10514 3238 10526 3290
rect 10526 3238 10556 3290
rect 10580 3238 10590 3290
rect 10590 3238 10636 3290
rect 10340 3236 10396 3238
rect 10420 3236 10476 3238
rect 10500 3236 10556 3238
rect 10580 3236 10636 3238
rect 8776 2746 8832 2748
rect 8856 2746 8912 2748
rect 8936 2746 8992 2748
rect 9016 2746 9072 2748
rect 8776 2694 8822 2746
rect 8822 2694 8832 2746
rect 8856 2694 8886 2746
rect 8886 2694 8898 2746
rect 8898 2694 8912 2746
rect 8936 2694 8950 2746
rect 8950 2694 8962 2746
rect 8962 2694 8992 2746
rect 9016 2694 9026 2746
rect 9026 2694 9072 2746
rect 8776 2692 8832 2694
rect 8856 2692 8912 2694
rect 8936 2692 8992 2694
rect 9016 2692 9072 2694
rect 11904 4922 11960 4924
rect 11984 4922 12040 4924
rect 12064 4922 12120 4924
rect 12144 4922 12200 4924
rect 11904 4870 11950 4922
rect 11950 4870 11960 4922
rect 11984 4870 12014 4922
rect 12014 4870 12026 4922
rect 12026 4870 12040 4922
rect 12064 4870 12078 4922
rect 12078 4870 12090 4922
rect 12090 4870 12120 4922
rect 12144 4870 12154 4922
rect 12154 4870 12200 4922
rect 11904 4868 11960 4870
rect 11984 4868 12040 4870
rect 12064 4868 12120 4870
rect 12144 4868 12200 4870
rect 12898 4800 12954 4856
rect 11904 3834 11960 3836
rect 11984 3834 12040 3836
rect 12064 3834 12120 3836
rect 12144 3834 12200 3836
rect 11904 3782 11950 3834
rect 11950 3782 11960 3834
rect 11984 3782 12014 3834
rect 12014 3782 12026 3834
rect 12026 3782 12040 3834
rect 12064 3782 12078 3834
rect 12078 3782 12090 3834
rect 12090 3782 12120 3834
rect 12144 3782 12154 3834
rect 12154 3782 12200 3834
rect 11904 3780 11960 3782
rect 11984 3780 12040 3782
rect 12064 3780 12120 3782
rect 12144 3780 12200 3782
rect 11904 2746 11960 2748
rect 11984 2746 12040 2748
rect 12064 2746 12120 2748
rect 12144 2746 12200 2748
rect 11904 2694 11950 2746
rect 11950 2694 11960 2746
rect 11984 2694 12014 2746
rect 12014 2694 12026 2746
rect 12026 2694 12040 2746
rect 12064 2694 12078 2746
rect 12078 2694 12090 2746
rect 12090 2694 12120 2746
rect 12144 2694 12154 2746
rect 12154 2694 12200 2746
rect 11904 2692 11960 2694
rect 11984 2692 12040 2694
rect 12064 2692 12120 2694
rect 12144 2692 12200 2694
rect 4084 2202 4140 2204
rect 4164 2202 4220 2204
rect 4244 2202 4300 2204
rect 4324 2202 4380 2204
rect 4084 2150 4130 2202
rect 4130 2150 4140 2202
rect 4164 2150 4194 2202
rect 4194 2150 4206 2202
rect 4206 2150 4220 2202
rect 4244 2150 4258 2202
rect 4258 2150 4270 2202
rect 4270 2150 4300 2202
rect 4324 2150 4334 2202
rect 4334 2150 4380 2202
rect 4084 2148 4140 2150
rect 4164 2148 4220 2150
rect 4244 2148 4300 2150
rect 4324 2148 4380 2150
rect 7212 2202 7268 2204
rect 7292 2202 7348 2204
rect 7372 2202 7428 2204
rect 7452 2202 7508 2204
rect 7212 2150 7258 2202
rect 7258 2150 7268 2202
rect 7292 2150 7322 2202
rect 7322 2150 7334 2202
rect 7334 2150 7348 2202
rect 7372 2150 7386 2202
rect 7386 2150 7398 2202
rect 7398 2150 7428 2202
rect 7452 2150 7462 2202
rect 7462 2150 7508 2202
rect 7212 2148 7268 2150
rect 7292 2148 7348 2150
rect 7372 2148 7428 2150
rect 7452 2148 7508 2150
rect 10340 2202 10396 2204
rect 10420 2202 10476 2204
rect 10500 2202 10556 2204
rect 10580 2202 10636 2204
rect 10340 2150 10386 2202
rect 10386 2150 10396 2202
rect 10420 2150 10450 2202
rect 10450 2150 10462 2202
rect 10462 2150 10476 2202
rect 10500 2150 10514 2202
rect 10514 2150 10526 2202
rect 10526 2150 10556 2202
rect 10580 2150 10590 2202
rect 10590 2150 10636 2202
rect 10340 2148 10396 2150
rect 10420 2148 10476 2150
rect 10500 2148 10556 2150
rect 10580 2148 10636 2150
rect 12346 720 12402 776
<< metal3 >>
rect 0 15738 800 15768
rect 1485 15738 1551 15741
rect 0 15736 1551 15738
rect 0 15680 1490 15736
rect 1546 15680 1551 15736
rect 0 15678 1551 15680
rect 0 15648 800 15678
rect 1485 15675 1551 15678
rect 2508 14720 2828 14721
rect 2508 14656 2516 14720
rect 2580 14656 2596 14720
rect 2660 14656 2676 14720
rect 2740 14656 2756 14720
rect 2820 14656 2828 14720
rect 2508 14655 2828 14656
rect 5636 14720 5956 14721
rect 5636 14656 5644 14720
rect 5708 14656 5724 14720
rect 5788 14656 5804 14720
rect 5868 14656 5884 14720
rect 5948 14656 5956 14720
rect 5636 14655 5956 14656
rect 8764 14720 9084 14721
rect 8764 14656 8772 14720
rect 8836 14656 8852 14720
rect 8916 14656 8932 14720
rect 8996 14656 9012 14720
rect 9076 14656 9084 14720
rect 8764 14655 9084 14656
rect 11892 14720 12212 14721
rect 11892 14656 11900 14720
rect 11964 14656 11980 14720
rect 12044 14656 12060 14720
rect 12124 14656 12140 14720
rect 12204 14656 12212 14720
rect 11892 14655 12212 14656
rect 4072 14176 4392 14177
rect 4072 14112 4080 14176
rect 4144 14112 4160 14176
rect 4224 14112 4240 14176
rect 4304 14112 4320 14176
rect 4384 14112 4392 14176
rect 4072 14111 4392 14112
rect 7200 14176 7520 14177
rect 7200 14112 7208 14176
rect 7272 14112 7288 14176
rect 7352 14112 7368 14176
rect 7432 14112 7448 14176
rect 7512 14112 7520 14176
rect 7200 14111 7520 14112
rect 10328 14176 10648 14177
rect 10328 14112 10336 14176
rect 10400 14112 10416 14176
rect 10480 14112 10496 14176
rect 10560 14112 10576 14176
rect 10640 14112 10648 14176
rect 10328 14111 10648 14112
rect 2508 13632 2828 13633
rect 2508 13568 2516 13632
rect 2580 13568 2596 13632
rect 2660 13568 2676 13632
rect 2740 13568 2756 13632
rect 2820 13568 2828 13632
rect 2508 13567 2828 13568
rect 5636 13632 5956 13633
rect 5636 13568 5644 13632
rect 5708 13568 5724 13632
rect 5788 13568 5804 13632
rect 5868 13568 5884 13632
rect 5948 13568 5956 13632
rect 5636 13567 5956 13568
rect 8764 13632 9084 13633
rect 8764 13568 8772 13632
rect 8836 13568 8852 13632
rect 8916 13568 8932 13632
rect 8996 13568 9012 13632
rect 9076 13568 9084 13632
rect 8764 13567 9084 13568
rect 11892 13632 12212 13633
rect 11892 13568 11900 13632
rect 11964 13568 11980 13632
rect 12044 13568 12060 13632
rect 12124 13568 12140 13632
rect 12204 13568 12212 13632
rect 11892 13567 12212 13568
rect 4072 13088 4392 13089
rect 4072 13024 4080 13088
rect 4144 13024 4160 13088
rect 4224 13024 4240 13088
rect 4304 13024 4320 13088
rect 4384 13024 4392 13088
rect 4072 13023 4392 13024
rect 7200 13088 7520 13089
rect 7200 13024 7208 13088
rect 7272 13024 7288 13088
rect 7352 13024 7368 13088
rect 7432 13024 7448 13088
rect 7512 13024 7520 13088
rect 7200 13023 7520 13024
rect 10328 13088 10648 13089
rect 10328 13024 10336 13088
rect 10400 13024 10416 13088
rect 10480 13024 10496 13088
rect 10560 13024 10576 13088
rect 10640 13024 10648 13088
rect 10328 13023 10648 13024
rect 12801 13018 12867 13021
rect 13944 13018 14744 13048
rect 12801 13016 14744 13018
rect 12801 12960 12806 13016
rect 12862 12960 14744 13016
rect 12801 12958 14744 12960
rect 12801 12955 12867 12958
rect 13944 12928 14744 12958
rect 2508 12544 2828 12545
rect 2508 12480 2516 12544
rect 2580 12480 2596 12544
rect 2660 12480 2676 12544
rect 2740 12480 2756 12544
rect 2820 12480 2828 12544
rect 2508 12479 2828 12480
rect 5636 12544 5956 12545
rect 5636 12480 5644 12544
rect 5708 12480 5724 12544
rect 5788 12480 5804 12544
rect 5868 12480 5884 12544
rect 5948 12480 5956 12544
rect 5636 12479 5956 12480
rect 8764 12544 9084 12545
rect 8764 12480 8772 12544
rect 8836 12480 8852 12544
rect 8916 12480 8932 12544
rect 8996 12480 9012 12544
rect 9076 12480 9084 12544
rect 8764 12479 9084 12480
rect 11892 12544 12212 12545
rect 11892 12480 11900 12544
rect 11964 12480 11980 12544
rect 12044 12480 12060 12544
rect 12124 12480 12140 12544
rect 12204 12480 12212 12544
rect 11892 12479 12212 12480
rect 4072 12000 4392 12001
rect 4072 11936 4080 12000
rect 4144 11936 4160 12000
rect 4224 11936 4240 12000
rect 4304 11936 4320 12000
rect 4384 11936 4392 12000
rect 4072 11935 4392 11936
rect 7200 12000 7520 12001
rect 7200 11936 7208 12000
rect 7272 11936 7288 12000
rect 7352 11936 7368 12000
rect 7432 11936 7448 12000
rect 7512 11936 7520 12000
rect 7200 11935 7520 11936
rect 10328 12000 10648 12001
rect 10328 11936 10336 12000
rect 10400 11936 10416 12000
rect 10480 11936 10496 12000
rect 10560 11936 10576 12000
rect 10640 11936 10648 12000
rect 10328 11935 10648 11936
rect 0 11658 800 11688
rect 1485 11658 1551 11661
rect 0 11656 1551 11658
rect 0 11600 1490 11656
rect 1546 11600 1551 11656
rect 0 11598 1551 11600
rect 0 11568 800 11598
rect 1485 11595 1551 11598
rect 2508 11456 2828 11457
rect 2508 11392 2516 11456
rect 2580 11392 2596 11456
rect 2660 11392 2676 11456
rect 2740 11392 2756 11456
rect 2820 11392 2828 11456
rect 2508 11391 2828 11392
rect 5636 11456 5956 11457
rect 5636 11392 5644 11456
rect 5708 11392 5724 11456
rect 5788 11392 5804 11456
rect 5868 11392 5884 11456
rect 5948 11392 5956 11456
rect 5636 11391 5956 11392
rect 8764 11456 9084 11457
rect 8764 11392 8772 11456
rect 8836 11392 8852 11456
rect 8916 11392 8932 11456
rect 8996 11392 9012 11456
rect 9076 11392 9084 11456
rect 8764 11391 9084 11392
rect 11892 11456 12212 11457
rect 11892 11392 11900 11456
rect 11964 11392 11980 11456
rect 12044 11392 12060 11456
rect 12124 11392 12140 11456
rect 12204 11392 12212 11456
rect 11892 11391 12212 11392
rect 4072 10912 4392 10913
rect 4072 10848 4080 10912
rect 4144 10848 4160 10912
rect 4224 10848 4240 10912
rect 4304 10848 4320 10912
rect 4384 10848 4392 10912
rect 4072 10847 4392 10848
rect 7200 10912 7520 10913
rect 7200 10848 7208 10912
rect 7272 10848 7288 10912
rect 7352 10848 7368 10912
rect 7432 10848 7448 10912
rect 7512 10848 7520 10912
rect 7200 10847 7520 10848
rect 10328 10912 10648 10913
rect 10328 10848 10336 10912
rect 10400 10848 10416 10912
rect 10480 10848 10496 10912
rect 10560 10848 10576 10912
rect 10640 10848 10648 10912
rect 10328 10847 10648 10848
rect 2508 10368 2828 10369
rect 2508 10304 2516 10368
rect 2580 10304 2596 10368
rect 2660 10304 2676 10368
rect 2740 10304 2756 10368
rect 2820 10304 2828 10368
rect 2508 10303 2828 10304
rect 5636 10368 5956 10369
rect 5636 10304 5644 10368
rect 5708 10304 5724 10368
rect 5788 10304 5804 10368
rect 5868 10304 5884 10368
rect 5948 10304 5956 10368
rect 5636 10303 5956 10304
rect 8764 10368 9084 10369
rect 8764 10304 8772 10368
rect 8836 10304 8852 10368
rect 8916 10304 8932 10368
rect 8996 10304 9012 10368
rect 9076 10304 9084 10368
rect 8764 10303 9084 10304
rect 11892 10368 12212 10369
rect 11892 10304 11900 10368
rect 11964 10304 11980 10368
rect 12044 10304 12060 10368
rect 12124 10304 12140 10368
rect 12204 10304 12212 10368
rect 11892 10303 12212 10304
rect 4072 9824 4392 9825
rect 4072 9760 4080 9824
rect 4144 9760 4160 9824
rect 4224 9760 4240 9824
rect 4304 9760 4320 9824
rect 4384 9760 4392 9824
rect 4072 9759 4392 9760
rect 7200 9824 7520 9825
rect 7200 9760 7208 9824
rect 7272 9760 7288 9824
rect 7352 9760 7368 9824
rect 7432 9760 7448 9824
rect 7512 9760 7520 9824
rect 7200 9759 7520 9760
rect 10328 9824 10648 9825
rect 10328 9760 10336 9824
rect 10400 9760 10416 9824
rect 10480 9760 10496 9824
rect 10560 9760 10576 9824
rect 10640 9760 10648 9824
rect 10328 9759 10648 9760
rect 2508 9280 2828 9281
rect 2508 9216 2516 9280
rect 2580 9216 2596 9280
rect 2660 9216 2676 9280
rect 2740 9216 2756 9280
rect 2820 9216 2828 9280
rect 2508 9215 2828 9216
rect 5636 9280 5956 9281
rect 5636 9216 5644 9280
rect 5708 9216 5724 9280
rect 5788 9216 5804 9280
rect 5868 9216 5884 9280
rect 5948 9216 5956 9280
rect 5636 9215 5956 9216
rect 8764 9280 9084 9281
rect 8764 9216 8772 9280
rect 8836 9216 8852 9280
rect 8916 9216 8932 9280
rect 8996 9216 9012 9280
rect 9076 9216 9084 9280
rect 8764 9215 9084 9216
rect 11892 9280 12212 9281
rect 11892 9216 11900 9280
rect 11964 9216 11980 9280
rect 12044 9216 12060 9280
rect 12124 9216 12140 9280
rect 12204 9216 12212 9280
rect 11892 9215 12212 9216
rect 12801 8938 12867 8941
rect 13944 8938 14744 8968
rect 12801 8936 14744 8938
rect 12801 8880 12806 8936
rect 12862 8880 14744 8936
rect 12801 8878 14744 8880
rect 12801 8875 12867 8878
rect 13944 8848 14744 8878
rect 4072 8736 4392 8737
rect 4072 8672 4080 8736
rect 4144 8672 4160 8736
rect 4224 8672 4240 8736
rect 4304 8672 4320 8736
rect 4384 8672 4392 8736
rect 4072 8671 4392 8672
rect 7200 8736 7520 8737
rect 7200 8672 7208 8736
rect 7272 8672 7288 8736
rect 7352 8672 7368 8736
rect 7432 8672 7448 8736
rect 7512 8672 7520 8736
rect 7200 8671 7520 8672
rect 10328 8736 10648 8737
rect 10328 8672 10336 8736
rect 10400 8672 10416 8736
rect 10480 8672 10496 8736
rect 10560 8672 10576 8736
rect 10640 8672 10648 8736
rect 10328 8671 10648 8672
rect 2508 8192 2828 8193
rect 2508 8128 2516 8192
rect 2580 8128 2596 8192
rect 2660 8128 2676 8192
rect 2740 8128 2756 8192
rect 2820 8128 2828 8192
rect 2508 8127 2828 8128
rect 5636 8192 5956 8193
rect 5636 8128 5644 8192
rect 5708 8128 5724 8192
rect 5788 8128 5804 8192
rect 5868 8128 5884 8192
rect 5948 8128 5956 8192
rect 5636 8127 5956 8128
rect 8764 8192 9084 8193
rect 8764 8128 8772 8192
rect 8836 8128 8852 8192
rect 8916 8128 8932 8192
rect 8996 8128 9012 8192
rect 9076 8128 9084 8192
rect 8764 8127 9084 8128
rect 11892 8192 12212 8193
rect 11892 8128 11900 8192
rect 11964 8128 11980 8192
rect 12044 8128 12060 8192
rect 12124 8128 12140 8192
rect 12204 8128 12212 8192
rect 11892 8127 12212 8128
rect 4072 7648 4392 7649
rect 0 7578 800 7608
rect 4072 7584 4080 7648
rect 4144 7584 4160 7648
rect 4224 7584 4240 7648
rect 4304 7584 4320 7648
rect 4384 7584 4392 7648
rect 4072 7583 4392 7584
rect 7200 7648 7520 7649
rect 7200 7584 7208 7648
rect 7272 7584 7288 7648
rect 7352 7584 7368 7648
rect 7432 7584 7448 7648
rect 7512 7584 7520 7648
rect 7200 7583 7520 7584
rect 10328 7648 10648 7649
rect 10328 7584 10336 7648
rect 10400 7584 10416 7648
rect 10480 7584 10496 7648
rect 10560 7584 10576 7648
rect 10640 7584 10648 7648
rect 10328 7583 10648 7584
rect 1485 7578 1551 7581
rect 0 7576 1551 7578
rect 0 7520 1490 7576
rect 1546 7520 1551 7576
rect 0 7518 1551 7520
rect 0 7488 800 7518
rect 1485 7515 1551 7518
rect 2508 7104 2828 7105
rect 2508 7040 2516 7104
rect 2580 7040 2596 7104
rect 2660 7040 2676 7104
rect 2740 7040 2756 7104
rect 2820 7040 2828 7104
rect 2508 7039 2828 7040
rect 5636 7104 5956 7105
rect 5636 7040 5644 7104
rect 5708 7040 5724 7104
rect 5788 7040 5804 7104
rect 5868 7040 5884 7104
rect 5948 7040 5956 7104
rect 5636 7039 5956 7040
rect 8764 7104 9084 7105
rect 8764 7040 8772 7104
rect 8836 7040 8852 7104
rect 8916 7040 8932 7104
rect 8996 7040 9012 7104
rect 9076 7040 9084 7104
rect 8764 7039 9084 7040
rect 11892 7104 12212 7105
rect 11892 7040 11900 7104
rect 11964 7040 11980 7104
rect 12044 7040 12060 7104
rect 12124 7040 12140 7104
rect 12204 7040 12212 7104
rect 11892 7039 12212 7040
rect 4072 6560 4392 6561
rect 4072 6496 4080 6560
rect 4144 6496 4160 6560
rect 4224 6496 4240 6560
rect 4304 6496 4320 6560
rect 4384 6496 4392 6560
rect 4072 6495 4392 6496
rect 7200 6560 7520 6561
rect 7200 6496 7208 6560
rect 7272 6496 7288 6560
rect 7352 6496 7368 6560
rect 7432 6496 7448 6560
rect 7512 6496 7520 6560
rect 7200 6495 7520 6496
rect 10328 6560 10648 6561
rect 10328 6496 10336 6560
rect 10400 6496 10416 6560
rect 10480 6496 10496 6560
rect 10560 6496 10576 6560
rect 10640 6496 10648 6560
rect 10328 6495 10648 6496
rect 2508 6016 2828 6017
rect 2508 5952 2516 6016
rect 2580 5952 2596 6016
rect 2660 5952 2676 6016
rect 2740 5952 2756 6016
rect 2820 5952 2828 6016
rect 2508 5951 2828 5952
rect 5636 6016 5956 6017
rect 5636 5952 5644 6016
rect 5708 5952 5724 6016
rect 5788 5952 5804 6016
rect 5868 5952 5884 6016
rect 5948 5952 5956 6016
rect 5636 5951 5956 5952
rect 8764 6016 9084 6017
rect 8764 5952 8772 6016
rect 8836 5952 8852 6016
rect 8916 5952 8932 6016
rect 8996 5952 9012 6016
rect 9076 5952 9084 6016
rect 8764 5951 9084 5952
rect 11892 6016 12212 6017
rect 11892 5952 11900 6016
rect 11964 5952 11980 6016
rect 12044 5952 12060 6016
rect 12124 5952 12140 6016
rect 12204 5952 12212 6016
rect 11892 5951 12212 5952
rect 4072 5472 4392 5473
rect 4072 5408 4080 5472
rect 4144 5408 4160 5472
rect 4224 5408 4240 5472
rect 4304 5408 4320 5472
rect 4384 5408 4392 5472
rect 4072 5407 4392 5408
rect 7200 5472 7520 5473
rect 7200 5408 7208 5472
rect 7272 5408 7288 5472
rect 7352 5408 7368 5472
rect 7432 5408 7448 5472
rect 7512 5408 7520 5472
rect 7200 5407 7520 5408
rect 10328 5472 10648 5473
rect 10328 5408 10336 5472
rect 10400 5408 10416 5472
rect 10480 5408 10496 5472
rect 10560 5408 10576 5472
rect 10640 5408 10648 5472
rect 10328 5407 10648 5408
rect 2508 4928 2828 4929
rect 2508 4864 2516 4928
rect 2580 4864 2596 4928
rect 2660 4864 2676 4928
rect 2740 4864 2756 4928
rect 2820 4864 2828 4928
rect 2508 4863 2828 4864
rect 5636 4928 5956 4929
rect 5636 4864 5644 4928
rect 5708 4864 5724 4928
rect 5788 4864 5804 4928
rect 5868 4864 5884 4928
rect 5948 4864 5956 4928
rect 5636 4863 5956 4864
rect 8764 4928 9084 4929
rect 8764 4864 8772 4928
rect 8836 4864 8852 4928
rect 8916 4864 8932 4928
rect 8996 4864 9012 4928
rect 9076 4864 9084 4928
rect 8764 4863 9084 4864
rect 11892 4928 12212 4929
rect 11892 4864 11900 4928
rect 11964 4864 11980 4928
rect 12044 4864 12060 4928
rect 12124 4864 12140 4928
rect 12204 4864 12212 4928
rect 11892 4863 12212 4864
rect 12893 4858 12959 4861
rect 13944 4858 14744 4888
rect 12893 4856 14744 4858
rect 12893 4800 12898 4856
rect 12954 4800 14744 4856
rect 12893 4798 14744 4800
rect 12893 4795 12959 4798
rect 13944 4768 14744 4798
rect 4072 4384 4392 4385
rect 4072 4320 4080 4384
rect 4144 4320 4160 4384
rect 4224 4320 4240 4384
rect 4304 4320 4320 4384
rect 4384 4320 4392 4384
rect 4072 4319 4392 4320
rect 7200 4384 7520 4385
rect 7200 4320 7208 4384
rect 7272 4320 7288 4384
rect 7352 4320 7368 4384
rect 7432 4320 7448 4384
rect 7512 4320 7520 4384
rect 7200 4319 7520 4320
rect 10328 4384 10648 4385
rect 10328 4320 10336 4384
rect 10400 4320 10416 4384
rect 10480 4320 10496 4384
rect 10560 4320 10576 4384
rect 10640 4320 10648 4384
rect 10328 4319 10648 4320
rect 2508 3840 2828 3841
rect 2508 3776 2516 3840
rect 2580 3776 2596 3840
rect 2660 3776 2676 3840
rect 2740 3776 2756 3840
rect 2820 3776 2828 3840
rect 2508 3775 2828 3776
rect 5636 3840 5956 3841
rect 5636 3776 5644 3840
rect 5708 3776 5724 3840
rect 5788 3776 5804 3840
rect 5868 3776 5884 3840
rect 5948 3776 5956 3840
rect 5636 3775 5956 3776
rect 8764 3840 9084 3841
rect 8764 3776 8772 3840
rect 8836 3776 8852 3840
rect 8916 3776 8932 3840
rect 8996 3776 9012 3840
rect 9076 3776 9084 3840
rect 8764 3775 9084 3776
rect 11892 3840 12212 3841
rect 11892 3776 11900 3840
rect 11964 3776 11980 3840
rect 12044 3776 12060 3840
rect 12124 3776 12140 3840
rect 12204 3776 12212 3840
rect 11892 3775 12212 3776
rect 0 3498 800 3528
rect 1485 3498 1551 3501
rect 0 3496 1551 3498
rect 0 3440 1490 3496
rect 1546 3440 1551 3496
rect 0 3438 1551 3440
rect 0 3408 800 3438
rect 1485 3435 1551 3438
rect 4072 3296 4392 3297
rect 4072 3232 4080 3296
rect 4144 3232 4160 3296
rect 4224 3232 4240 3296
rect 4304 3232 4320 3296
rect 4384 3232 4392 3296
rect 4072 3231 4392 3232
rect 7200 3296 7520 3297
rect 7200 3232 7208 3296
rect 7272 3232 7288 3296
rect 7352 3232 7368 3296
rect 7432 3232 7448 3296
rect 7512 3232 7520 3296
rect 7200 3231 7520 3232
rect 10328 3296 10648 3297
rect 10328 3232 10336 3296
rect 10400 3232 10416 3296
rect 10480 3232 10496 3296
rect 10560 3232 10576 3296
rect 10640 3232 10648 3296
rect 10328 3231 10648 3232
rect 2508 2752 2828 2753
rect 2508 2688 2516 2752
rect 2580 2688 2596 2752
rect 2660 2688 2676 2752
rect 2740 2688 2756 2752
rect 2820 2688 2828 2752
rect 2508 2687 2828 2688
rect 5636 2752 5956 2753
rect 5636 2688 5644 2752
rect 5708 2688 5724 2752
rect 5788 2688 5804 2752
rect 5868 2688 5884 2752
rect 5948 2688 5956 2752
rect 5636 2687 5956 2688
rect 8764 2752 9084 2753
rect 8764 2688 8772 2752
rect 8836 2688 8852 2752
rect 8916 2688 8932 2752
rect 8996 2688 9012 2752
rect 9076 2688 9084 2752
rect 8764 2687 9084 2688
rect 11892 2752 12212 2753
rect 11892 2688 11900 2752
rect 11964 2688 11980 2752
rect 12044 2688 12060 2752
rect 12124 2688 12140 2752
rect 12204 2688 12212 2752
rect 11892 2687 12212 2688
rect 4072 2208 4392 2209
rect 4072 2144 4080 2208
rect 4144 2144 4160 2208
rect 4224 2144 4240 2208
rect 4304 2144 4320 2208
rect 4384 2144 4392 2208
rect 4072 2143 4392 2144
rect 7200 2208 7520 2209
rect 7200 2144 7208 2208
rect 7272 2144 7288 2208
rect 7352 2144 7368 2208
rect 7432 2144 7448 2208
rect 7512 2144 7520 2208
rect 7200 2143 7520 2144
rect 10328 2208 10648 2209
rect 10328 2144 10336 2208
rect 10400 2144 10416 2208
rect 10480 2144 10496 2208
rect 10560 2144 10576 2208
rect 10640 2144 10648 2208
rect 10328 2143 10648 2144
rect 12341 778 12407 781
rect 13944 778 14744 808
rect 12341 776 14744 778
rect 12341 720 12346 776
rect 12402 720 14744 776
rect 12341 718 14744 720
rect 12341 715 12407 718
rect 13944 688 14744 718
<< via3 >>
rect 2516 14716 2580 14720
rect 2516 14660 2520 14716
rect 2520 14660 2576 14716
rect 2576 14660 2580 14716
rect 2516 14656 2580 14660
rect 2596 14716 2660 14720
rect 2596 14660 2600 14716
rect 2600 14660 2656 14716
rect 2656 14660 2660 14716
rect 2596 14656 2660 14660
rect 2676 14716 2740 14720
rect 2676 14660 2680 14716
rect 2680 14660 2736 14716
rect 2736 14660 2740 14716
rect 2676 14656 2740 14660
rect 2756 14716 2820 14720
rect 2756 14660 2760 14716
rect 2760 14660 2816 14716
rect 2816 14660 2820 14716
rect 2756 14656 2820 14660
rect 5644 14716 5708 14720
rect 5644 14660 5648 14716
rect 5648 14660 5704 14716
rect 5704 14660 5708 14716
rect 5644 14656 5708 14660
rect 5724 14716 5788 14720
rect 5724 14660 5728 14716
rect 5728 14660 5784 14716
rect 5784 14660 5788 14716
rect 5724 14656 5788 14660
rect 5804 14716 5868 14720
rect 5804 14660 5808 14716
rect 5808 14660 5864 14716
rect 5864 14660 5868 14716
rect 5804 14656 5868 14660
rect 5884 14716 5948 14720
rect 5884 14660 5888 14716
rect 5888 14660 5944 14716
rect 5944 14660 5948 14716
rect 5884 14656 5948 14660
rect 8772 14716 8836 14720
rect 8772 14660 8776 14716
rect 8776 14660 8832 14716
rect 8832 14660 8836 14716
rect 8772 14656 8836 14660
rect 8852 14716 8916 14720
rect 8852 14660 8856 14716
rect 8856 14660 8912 14716
rect 8912 14660 8916 14716
rect 8852 14656 8916 14660
rect 8932 14716 8996 14720
rect 8932 14660 8936 14716
rect 8936 14660 8992 14716
rect 8992 14660 8996 14716
rect 8932 14656 8996 14660
rect 9012 14716 9076 14720
rect 9012 14660 9016 14716
rect 9016 14660 9072 14716
rect 9072 14660 9076 14716
rect 9012 14656 9076 14660
rect 11900 14716 11964 14720
rect 11900 14660 11904 14716
rect 11904 14660 11960 14716
rect 11960 14660 11964 14716
rect 11900 14656 11964 14660
rect 11980 14716 12044 14720
rect 11980 14660 11984 14716
rect 11984 14660 12040 14716
rect 12040 14660 12044 14716
rect 11980 14656 12044 14660
rect 12060 14716 12124 14720
rect 12060 14660 12064 14716
rect 12064 14660 12120 14716
rect 12120 14660 12124 14716
rect 12060 14656 12124 14660
rect 12140 14716 12204 14720
rect 12140 14660 12144 14716
rect 12144 14660 12200 14716
rect 12200 14660 12204 14716
rect 12140 14656 12204 14660
rect 4080 14172 4144 14176
rect 4080 14116 4084 14172
rect 4084 14116 4140 14172
rect 4140 14116 4144 14172
rect 4080 14112 4144 14116
rect 4160 14172 4224 14176
rect 4160 14116 4164 14172
rect 4164 14116 4220 14172
rect 4220 14116 4224 14172
rect 4160 14112 4224 14116
rect 4240 14172 4304 14176
rect 4240 14116 4244 14172
rect 4244 14116 4300 14172
rect 4300 14116 4304 14172
rect 4240 14112 4304 14116
rect 4320 14172 4384 14176
rect 4320 14116 4324 14172
rect 4324 14116 4380 14172
rect 4380 14116 4384 14172
rect 4320 14112 4384 14116
rect 7208 14172 7272 14176
rect 7208 14116 7212 14172
rect 7212 14116 7268 14172
rect 7268 14116 7272 14172
rect 7208 14112 7272 14116
rect 7288 14172 7352 14176
rect 7288 14116 7292 14172
rect 7292 14116 7348 14172
rect 7348 14116 7352 14172
rect 7288 14112 7352 14116
rect 7368 14172 7432 14176
rect 7368 14116 7372 14172
rect 7372 14116 7428 14172
rect 7428 14116 7432 14172
rect 7368 14112 7432 14116
rect 7448 14172 7512 14176
rect 7448 14116 7452 14172
rect 7452 14116 7508 14172
rect 7508 14116 7512 14172
rect 7448 14112 7512 14116
rect 10336 14172 10400 14176
rect 10336 14116 10340 14172
rect 10340 14116 10396 14172
rect 10396 14116 10400 14172
rect 10336 14112 10400 14116
rect 10416 14172 10480 14176
rect 10416 14116 10420 14172
rect 10420 14116 10476 14172
rect 10476 14116 10480 14172
rect 10416 14112 10480 14116
rect 10496 14172 10560 14176
rect 10496 14116 10500 14172
rect 10500 14116 10556 14172
rect 10556 14116 10560 14172
rect 10496 14112 10560 14116
rect 10576 14172 10640 14176
rect 10576 14116 10580 14172
rect 10580 14116 10636 14172
rect 10636 14116 10640 14172
rect 10576 14112 10640 14116
rect 2516 13628 2580 13632
rect 2516 13572 2520 13628
rect 2520 13572 2576 13628
rect 2576 13572 2580 13628
rect 2516 13568 2580 13572
rect 2596 13628 2660 13632
rect 2596 13572 2600 13628
rect 2600 13572 2656 13628
rect 2656 13572 2660 13628
rect 2596 13568 2660 13572
rect 2676 13628 2740 13632
rect 2676 13572 2680 13628
rect 2680 13572 2736 13628
rect 2736 13572 2740 13628
rect 2676 13568 2740 13572
rect 2756 13628 2820 13632
rect 2756 13572 2760 13628
rect 2760 13572 2816 13628
rect 2816 13572 2820 13628
rect 2756 13568 2820 13572
rect 5644 13628 5708 13632
rect 5644 13572 5648 13628
rect 5648 13572 5704 13628
rect 5704 13572 5708 13628
rect 5644 13568 5708 13572
rect 5724 13628 5788 13632
rect 5724 13572 5728 13628
rect 5728 13572 5784 13628
rect 5784 13572 5788 13628
rect 5724 13568 5788 13572
rect 5804 13628 5868 13632
rect 5804 13572 5808 13628
rect 5808 13572 5864 13628
rect 5864 13572 5868 13628
rect 5804 13568 5868 13572
rect 5884 13628 5948 13632
rect 5884 13572 5888 13628
rect 5888 13572 5944 13628
rect 5944 13572 5948 13628
rect 5884 13568 5948 13572
rect 8772 13628 8836 13632
rect 8772 13572 8776 13628
rect 8776 13572 8832 13628
rect 8832 13572 8836 13628
rect 8772 13568 8836 13572
rect 8852 13628 8916 13632
rect 8852 13572 8856 13628
rect 8856 13572 8912 13628
rect 8912 13572 8916 13628
rect 8852 13568 8916 13572
rect 8932 13628 8996 13632
rect 8932 13572 8936 13628
rect 8936 13572 8992 13628
rect 8992 13572 8996 13628
rect 8932 13568 8996 13572
rect 9012 13628 9076 13632
rect 9012 13572 9016 13628
rect 9016 13572 9072 13628
rect 9072 13572 9076 13628
rect 9012 13568 9076 13572
rect 11900 13628 11964 13632
rect 11900 13572 11904 13628
rect 11904 13572 11960 13628
rect 11960 13572 11964 13628
rect 11900 13568 11964 13572
rect 11980 13628 12044 13632
rect 11980 13572 11984 13628
rect 11984 13572 12040 13628
rect 12040 13572 12044 13628
rect 11980 13568 12044 13572
rect 12060 13628 12124 13632
rect 12060 13572 12064 13628
rect 12064 13572 12120 13628
rect 12120 13572 12124 13628
rect 12060 13568 12124 13572
rect 12140 13628 12204 13632
rect 12140 13572 12144 13628
rect 12144 13572 12200 13628
rect 12200 13572 12204 13628
rect 12140 13568 12204 13572
rect 4080 13084 4144 13088
rect 4080 13028 4084 13084
rect 4084 13028 4140 13084
rect 4140 13028 4144 13084
rect 4080 13024 4144 13028
rect 4160 13084 4224 13088
rect 4160 13028 4164 13084
rect 4164 13028 4220 13084
rect 4220 13028 4224 13084
rect 4160 13024 4224 13028
rect 4240 13084 4304 13088
rect 4240 13028 4244 13084
rect 4244 13028 4300 13084
rect 4300 13028 4304 13084
rect 4240 13024 4304 13028
rect 4320 13084 4384 13088
rect 4320 13028 4324 13084
rect 4324 13028 4380 13084
rect 4380 13028 4384 13084
rect 4320 13024 4384 13028
rect 7208 13084 7272 13088
rect 7208 13028 7212 13084
rect 7212 13028 7268 13084
rect 7268 13028 7272 13084
rect 7208 13024 7272 13028
rect 7288 13084 7352 13088
rect 7288 13028 7292 13084
rect 7292 13028 7348 13084
rect 7348 13028 7352 13084
rect 7288 13024 7352 13028
rect 7368 13084 7432 13088
rect 7368 13028 7372 13084
rect 7372 13028 7428 13084
rect 7428 13028 7432 13084
rect 7368 13024 7432 13028
rect 7448 13084 7512 13088
rect 7448 13028 7452 13084
rect 7452 13028 7508 13084
rect 7508 13028 7512 13084
rect 7448 13024 7512 13028
rect 10336 13084 10400 13088
rect 10336 13028 10340 13084
rect 10340 13028 10396 13084
rect 10396 13028 10400 13084
rect 10336 13024 10400 13028
rect 10416 13084 10480 13088
rect 10416 13028 10420 13084
rect 10420 13028 10476 13084
rect 10476 13028 10480 13084
rect 10416 13024 10480 13028
rect 10496 13084 10560 13088
rect 10496 13028 10500 13084
rect 10500 13028 10556 13084
rect 10556 13028 10560 13084
rect 10496 13024 10560 13028
rect 10576 13084 10640 13088
rect 10576 13028 10580 13084
rect 10580 13028 10636 13084
rect 10636 13028 10640 13084
rect 10576 13024 10640 13028
rect 2516 12540 2580 12544
rect 2516 12484 2520 12540
rect 2520 12484 2576 12540
rect 2576 12484 2580 12540
rect 2516 12480 2580 12484
rect 2596 12540 2660 12544
rect 2596 12484 2600 12540
rect 2600 12484 2656 12540
rect 2656 12484 2660 12540
rect 2596 12480 2660 12484
rect 2676 12540 2740 12544
rect 2676 12484 2680 12540
rect 2680 12484 2736 12540
rect 2736 12484 2740 12540
rect 2676 12480 2740 12484
rect 2756 12540 2820 12544
rect 2756 12484 2760 12540
rect 2760 12484 2816 12540
rect 2816 12484 2820 12540
rect 2756 12480 2820 12484
rect 5644 12540 5708 12544
rect 5644 12484 5648 12540
rect 5648 12484 5704 12540
rect 5704 12484 5708 12540
rect 5644 12480 5708 12484
rect 5724 12540 5788 12544
rect 5724 12484 5728 12540
rect 5728 12484 5784 12540
rect 5784 12484 5788 12540
rect 5724 12480 5788 12484
rect 5804 12540 5868 12544
rect 5804 12484 5808 12540
rect 5808 12484 5864 12540
rect 5864 12484 5868 12540
rect 5804 12480 5868 12484
rect 5884 12540 5948 12544
rect 5884 12484 5888 12540
rect 5888 12484 5944 12540
rect 5944 12484 5948 12540
rect 5884 12480 5948 12484
rect 8772 12540 8836 12544
rect 8772 12484 8776 12540
rect 8776 12484 8832 12540
rect 8832 12484 8836 12540
rect 8772 12480 8836 12484
rect 8852 12540 8916 12544
rect 8852 12484 8856 12540
rect 8856 12484 8912 12540
rect 8912 12484 8916 12540
rect 8852 12480 8916 12484
rect 8932 12540 8996 12544
rect 8932 12484 8936 12540
rect 8936 12484 8992 12540
rect 8992 12484 8996 12540
rect 8932 12480 8996 12484
rect 9012 12540 9076 12544
rect 9012 12484 9016 12540
rect 9016 12484 9072 12540
rect 9072 12484 9076 12540
rect 9012 12480 9076 12484
rect 11900 12540 11964 12544
rect 11900 12484 11904 12540
rect 11904 12484 11960 12540
rect 11960 12484 11964 12540
rect 11900 12480 11964 12484
rect 11980 12540 12044 12544
rect 11980 12484 11984 12540
rect 11984 12484 12040 12540
rect 12040 12484 12044 12540
rect 11980 12480 12044 12484
rect 12060 12540 12124 12544
rect 12060 12484 12064 12540
rect 12064 12484 12120 12540
rect 12120 12484 12124 12540
rect 12060 12480 12124 12484
rect 12140 12540 12204 12544
rect 12140 12484 12144 12540
rect 12144 12484 12200 12540
rect 12200 12484 12204 12540
rect 12140 12480 12204 12484
rect 4080 11996 4144 12000
rect 4080 11940 4084 11996
rect 4084 11940 4140 11996
rect 4140 11940 4144 11996
rect 4080 11936 4144 11940
rect 4160 11996 4224 12000
rect 4160 11940 4164 11996
rect 4164 11940 4220 11996
rect 4220 11940 4224 11996
rect 4160 11936 4224 11940
rect 4240 11996 4304 12000
rect 4240 11940 4244 11996
rect 4244 11940 4300 11996
rect 4300 11940 4304 11996
rect 4240 11936 4304 11940
rect 4320 11996 4384 12000
rect 4320 11940 4324 11996
rect 4324 11940 4380 11996
rect 4380 11940 4384 11996
rect 4320 11936 4384 11940
rect 7208 11996 7272 12000
rect 7208 11940 7212 11996
rect 7212 11940 7268 11996
rect 7268 11940 7272 11996
rect 7208 11936 7272 11940
rect 7288 11996 7352 12000
rect 7288 11940 7292 11996
rect 7292 11940 7348 11996
rect 7348 11940 7352 11996
rect 7288 11936 7352 11940
rect 7368 11996 7432 12000
rect 7368 11940 7372 11996
rect 7372 11940 7428 11996
rect 7428 11940 7432 11996
rect 7368 11936 7432 11940
rect 7448 11996 7512 12000
rect 7448 11940 7452 11996
rect 7452 11940 7508 11996
rect 7508 11940 7512 11996
rect 7448 11936 7512 11940
rect 10336 11996 10400 12000
rect 10336 11940 10340 11996
rect 10340 11940 10396 11996
rect 10396 11940 10400 11996
rect 10336 11936 10400 11940
rect 10416 11996 10480 12000
rect 10416 11940 10420 11996
rect 10420 11940 10476 11996
rect 10476 11940 10480 11996
rect 10416 11936 10480 11940
rect 10496 11996 10560 12000
rect 10496 11940 10500 11996
rect 10500 11940 10556 11996
rect 10556 11940 10560 11996
rect 10496 11936 10560 11940
rect 10576 11996 10640 12000
rect 10576 11940 10580 11996
rect 10580 11940 10636 11996
rect 10636 11940 10640 11996
rect 10576 11936 10640 11940
rect 2516 11452 2580 11456
rect 2516 11396 2520 11452
rect 2520 11396 2576 11452
rect 2576 11396 2580 11452
rect 2516 11392 2580 11396
rect 2596 11452 2660 11456
rect 2596 11396 2600 11452
rect 2600 11396 2656 11452
rect 2656 11396 2660 11452
rect 2596 11392 2660 11396
rect 2676 11452 2740 11456
rect 2676 11396 2680 11452
rect 2680 11396 2736 11452
rect 2736 11396 2740 11452
rect 2676 11392 2740 11396
rect 2756 11452 2820 11456
rect 2756 11396 2760 11452
rect 2760 11396 2816 11452
rect 2816 11396 2820 11452
rect 2756 11392 2820 11396
rect 5644 11452 5708 11456
rect 5644 11396 5648 11452
rect 5648 11396 5704 11452
rect 5704 11396 5708 11452
rect 5644 11392 5708 11396
rect 5724 11452 5788 11456
rect 5724 11396 5728 11452
rect 5728 11396 5784 11452
rect 5784 11396 5788 11452
rect 5724 11392 5788 11396
rect 5804 11452 5868 11456
rect 5804 11396 5808 11452
rect 5808 11396 5864 11452
rect 5864 11396 5868 11452
rect 5804 11392 5868 11396
rect 5884 11452 5948 11456
rect 5884 11396 5888 11452
rect 5888 11396 5944 11452
rect 5944 11396 5948 11452
rect 5884 11392 5948 11396
rect 8772 11452 8836 11456
rect 8772 11396 8776 11452
rect 8776 11396 8832 11452
rect 8832 11396 8836 11452
rect 8772 11392 8836 11396
rect 8852 11452 8916 11456
rect 8852 11396 8856 11452
rect 8856 11396 8912 11452
rect 8912 11396 8916 11452
rect 8852 11392 8916 11396
rect 8932 11452 8996 11456
rect 8932 11396 8936 11452
rect 8936 11396 8992 11452
rect 8992 11396 8996 11452
rect 8932 11392 8996 11396
rect 9012 11452 9076 11456
rect 9012 11396 9016 11452
rect 9016 11396 9072 11452
rect 9072 11396 9076 11452
rect 9012 11392 9076 11396
rect 11900 11452 11964 11456
rect 11900 11396 11904 11452
rect 11904 11396 11960 11452
rect 11960 11396 11964 11452
rect 11900 11392 11964 11396
rect 11980 11452 12044 11456
rect 11980 11396 11984 11452
rect 11984 11396 12040 11452
rect 12040 11396 12044 11452
rect 11980 11392 12044 11396
rect 12060 11452 12124 11456
rect 12060 11396 12064 11452
rect 12064 11396 12120 11452
rect 12120 11396 12124 11452
rect 12060 11392 12124 11396
rect 12140 11452 12204 11456
rect 12140 11396 12144 11452
rect 12144 11396 12200 11452
rect 12200 11396 12204 11452
rect 12140 11392 12204 11396
rect 4080 10908 4144 10912
rect 4080 10852 4084 10908
rect 4084 10852 4140 10908
rect 4140 10852 4144 10908
rect 4080 10848 4144 10852
rect 4160 10908 4224 10912
rect 4160 10852 4164 10908
rect 4164 10852 4220 10908
rect 4220 10852 4224 10908
rect 4160 10848 4224 10852
rect 4240 10908 4304 10912
rect 4240 10852 4244 10908
rect 4244 10852 4300 10908
rect 4300 10852 4304 10908
rect 4240 10848 4304 10852
rect 4320 10908 4384 10912
rect 4320 10852 4324 10908
rect 4324 10852 4380 10908
rect 4380 10852 4384 10908
rect 4320 10848 4384 10852
rect 7208 10908 7272 10912
rect 7208 10852 7212 10908
rect 7212 10852 7268 10908
rect 7268 10852 7272 10908
rect 7208 10848 7272 10852
rect 7288 10908 7352 10912
rect 7288 10852 7292 10908
rect 7292 10852 7348 10908
rect 7348 10852 7352 10908
rect 7288 10848 7352 10852
rect 7368 10908 7432 10912
rect 7368 10852 7372 10908
rect 7372 10852 7428 10908
rect 7428 10852 7432 10908
rect 7368 10848 7432 10852
rect 7448 10908 7512 10912
rect 7448 10852 7452 10908
rect 7452 10852 7508 10908
rect 7508 10852 7512 10908
rect 7448 10848 7512 10852
rect 10336 10908 10400 10912
rect 10336 10852 10340 10908
rect 10340 10852 10396 10908
rect 10396 10852 10400 10908
rect 10336 10848 10400 10852
rect 10416 10908 10480 10912
rect 10416 10852 10420 10908
rect 10420 10852 10476 10908
rect 10476 10852 10480 10908
rect 10416 10848 10480 10852
rect 10496 10908 10560 10912
rect 10496 10852 10500 10908
rect 10500 10852 10556 10908
rect 10556 10852 10560 10908
rect 10496 10848 10560 10852
rect 10576 10908 10640 10912
rect 10576 10852 10580 10908
rect 10580 10852 10636 10908
rect 10636 10852 10640 10908
rect 10576 10848 10640 10852
rect 2516 10364 2580 10368
rect 2516 10308 2520 10364
rect 2520 10308 2576 10364
rect 2576 10308 2580 10364
rect 2516 10304 2580 10308
rect 2596 10364 2660 10368
rect 2596 10308 2600 10364
rect 2600 10308 2656 10364
rect 2656 10308 2660 10364
rect 2596 10304 2660 10308
rect 2676 10364 2740 10368
rect 2676 10308 2680 10364
rect 2680 10308 2736 10364
rect 2736 10308 2740 10364
rect 2676 10304 2740 10308
rect 2756 10364 2820 10368
rect 2756 10308 2760 10364
rect 2760 10308 2816 10364
rect 2816 10308 2820 10364
rect 2756 10304 2820 10308
rect 5644 10364 5708 10368
rect 5644 10308 5648 10364
rect 5648 10308 5704 10364
rect 5704 10308 5708 10364
rect 5644 10304 5708 10308
rect 5724 10364 5788 10368
rect 5724 10308 5728 10364
rect 5728 10308 5784 10364
rect 5784 10308 5788 10364
rect 5724 10304 5788 10308
rect 5804 10364 5868 10368
rect 5804 10308 5808 10364
rect 5808 10308 5864 10364
rect 5864 10308 5868 10364
rect 5804 10304 5868 10308
rect 5884 10364 5948 10368
rect 5884 10308 5888 10364
rect 5888 10308 5944 10364
rect 5944 10308 5948 10364
rect 5884 10304 5948 10308
rect 8772 10364 8836 10368
rect 8772 10308 8776 10364
rect 8776 10308 8832 10364
rect 8832 10308 8836 10364
rect 8772 10304 8836 10308
rect 8852 10364 8916 10368
rect 8852 10308 8856 10364
rect 8856 10308 8912 10364
rect 8912 10308 8916 10364
rect 8852 10304 8916 10308
rect 8932 10364 8996 10368
rect 8932 10308 8936 10364
rect 8936 10308 8992 10364
rect 8992 10308 8996 10364
rect 8932 10304 8996 10308
rect 9012 10364 9076 10368
rect 9012 10308 9016 10364
rect 9016 10308 9072 10364
rect 9072 10308 9076 10364
rect 9012 10304 9076 10308
rect 11900 10364 11964 10368
rect 11900 10308 11904 10364
rect 11904 10308 11960 10364
rect 11960 10308 11964 10364
rect 11900 10304 11964 10308
rect 11980 10364 12044 10368
rect 11980 10308 11984 10364
rect 11984 10308 12040 10364
rect 12040 10308 12044 10364
rect 11980 10304 12044 10308
rect 12060 10364 12124 10368
rect 12060 10308 12064 10364
rect 12064 10308 12120 10364
rect 12120 10308 12124 10364
rect 12060 10304 12124 10308
rect 12140 10364 12204 10368
rect 12140 10308 12144 10364
rect 12144 10308 12200 10364
rect 12200 10308 12204 10364
rect 12140 10304 12204 10308
rect 4080 9820 4144 9824
rect 4080 9764 4084 9820
rect 4084 9764 4140 9820
rect 4140 9764 4144 9820
rect 4080 9760 4144 9764
rect 4160 9820 4224 9824
rect 4160 9764 4164 9820
rect 4164 9764 4220 9820
rect 4220 9764 4224 9820
rect 4160 9760 4224 9764
rect 4240 9820 4304 9824
rect 4240 9764 4244 9820
rect 4244 9764 4300 9820
rect 4300 9764 4304 9820
rect 4240 9760 4304 9764
rect 4320 9820 4384 9824
rect 4320 9764 4324 9820
rect 4324 9764 4380 9820
rect 4380 9764 4384 9820
rect 4320 9760 4384 9764
rect 7208 9820 7272 9824
rect 7208 9764 7212 9820
rect 7212 9764 7268 9820
rect 7268 9764 7272 9820
rect 7208 9760 7272 9764
rect 7288 9820 7352 9824
rect 7288 9764 7292 9820
rect 7292 9764 7348 9820
rect 7348 9764 7352 9820
rect 7288 9760 7352 9764
rect 7368 9820 7432 9824
rect 7368 9764 7372 9820
rect 7372 9764 7428 9820
rect 7428 9764 7432 9820
rect 7368 9760 7432 9764
rect 7448 9820 7512 9824
rect 7448 9764 7452 9820
rect 7452 9764 7508 9820
rect 7508 9764 7512 9820
rect 7448 9760 7512 9764
rect 10336 9820 10400 9824
rect 10336 9764 10340 9820
rect 10340 9764 10396 9820
rect 10396 9764 10400 9820
rect 10336 9760 10400 9764
rect 10416 9820 10480 9824
rect 10416 9764 10420 9820
rect 10420 9764 10476 9820
rect 10476 9764 10480 9820
rect 10416 9760 10480 9764
rect 10496 9820 10560 9824
rect 10496 9764 10500 9820
rect 10500 9764 10556 9820
rect 10556 9764 10560 9820
rect 10496 9760 10560 9764
rect 10576 9820 10640 9824
rect 10576 9764 10580 9820
rect 10580 9764 10636 9820
rect 10636 9764 10640 9820
rect 10576 9760 10640 9764
rect 2516 9276 2580 9280
rect 2516 9220 2520 9276
rect 2520 9220 2576 9276
rect 2576 9220 2580 9276
rect 2516 9216 2580 9220
rect 2596 9276 2660 9280
rect 2596 9220 2600 9276
rect 2600 9220 2656 9276
rect 2656 9220 2660 9276
rect 2596 9216 2660 9220
rect 2676 9276 2740 9280
rect 2676 9220 2680 9276
rect 2680 9220 2736 9276
rect 2736 9220 2740 9276
rect 2676 9216 2740 9220
rect 2756 9276 2820 9280
rect 2756 9220 2760 9276
rect 2760 9220 2816 9276
rect 2816 9220 2820 9276
rect 2756 9216 2820 9220
rect 5644 9276 5708 9280
rect 5644 9220 5648 9276
rect 5648 9220 5704 9276
rect 5704 9220 5708 9276
rect 5644 9216 5708 9220
rect 5724 9276 5788 9280
rect 5724 9220 5728 9276
rect 5728 9220 5784 9276
rect 5784 9220 5788 9276
rect 5724 9216 5788 9220
rect 5804 9276 5868 9280
rect 5804 9220 5808 9276
rect 5808 9220 5864 9276
rect 5864 9220 5868 9276
rect 5804 9216 5868 9220
rect 5884 9276 5948 9280
rect 5884 9220 5888 9276
rect 5888 9220 5944 9276
rect 5944 9220 5948 9276
rect 5884 9216 5948 9220
rect 8772 9276 8836 9280
rect 8772 9220 8776 9276
rect 8776 9220 8832 9276
rect 8832 9220 8836 9276
rect 8772 9216 8836 9220
rect 8852 9276 8916 9280
rect 8852 9220 8856 9276
rect 8856 9220 8912 9276
rect 8912 9220 8916 9276
rect 8852 9216 8916 9220
rect 8932 9276 8996 9280
rect 8932 9220 8936 9276
rect 8936 9220 8992 9276
rect 8992 9220 8996 9276
rect 8932 9216 8996 9220
rect 9012 9276 9076 9280
rect 9012 9220 9016 9276
rect 9016 9220 9072 9276
rect 9072 9220 9076 9276
rect 9012 9216 9076 9220
rect 11900 9276 11964 9280
rect 11900 9220 11904 9276
rect 11904 9220 11960 9276
rect 11960 9220 11964 9276
rect 11900 9216 11964 9220
rect 11980 9276 12044 9280
rect 11980 9220 11984 9276
rect 11984 9220 12040 9276
rect 12040 9220 12044 9276
rect 11980 9216 12044 9220
rect 12060 9276 12124 9280
rect 12060 9220 12064 9276
rect 12064 9220 12120 9276
rect 12120 9220 12124 9276
rect 12060 9216 12124 9220
rect 12140 9276 12204 9280
rect 12140 9220 12144 9276
rect 12144 9220 12200 9276
rect 12200 9220 12204 9276
rect 12140 9216 12204 9220
rect 4080 8732 4144 8736
rect 4080 8676 4084 8732
rect 4084 8676 4140 8732
rect 4140 8676 4144 8732
rect 4080 8672 4144 8676
rect 4160 8732 4224 8736
rect 4160 8676 4164 8732
rect 4164 8676 4220 8732
rect 4220 8676 4224 8732
rect 4160 8672 4224 8676
rect 4240 8732 4304 8736
rect 4240 8676 4244 8732
rect 4244 8676 4300 8732
rect 4300 8676 4304 8732
rect 4240 8672 4304 8676
rect 4320 8732 4384 8736
rect 4320 8676 4324 8732
rect 4324 8676 4380 8732
rect 4380 8676 4384 8732
rect 4320 8672 4384 8676
rect 7208 8732 7272 8736
rect 7208 8676 7212 8732
rect 7212 8676 7268 8732
rect 7268 8676 7272 8732
rect 7208 8672 7272 8676
rect 7288 8732 7352 8736
rect 7288 8676 7292 8732
rect 7292 8676 7348 8732
rect 7348 8676 7352 8732
rect 7288 8672 7352 8676
rect 7368 8732 7432 8736
rect 7368 8676 7372 8732
rect 7372 8676 7428 8732
rect 7428 8676 7432 8732
rect 7368 8672 7432 8676
rect 7448 8732 7512 8736
rect 7448 8676 7452 8732
rect 7452 8676 7508 8732
rect 7508 8676 7512 8732
rect 7448 8672 7512 8676
rect 10336 8732 10400 8736
rect 10336 8676 10340 8732
rect 10340 8676 10396 8732
rect 10396 8676 10400 8732
rect 10336 8672 10400 8676
rect 10416 8732 10480 8736
rect 10416 8676 10420 8732
rect 10420 8676 10476 8732
rect 10476 8676 10480 8732
rect 10416 8672 10480 8676
rect 10496 8732 10560 8736
rect 10496 8676 10500 8732
rect 10500 8676 10556 8732
rect 10556 8676 10560 8732
rect 10496 8672 10560 8676
rect 10576 8732 10640 8736
rect 10576 8676 10580 8732
rect 10580 8676 10636 8732
rect 10636 8676 10640 8732
rect 10576 8672 10640 8676
rect 2516 8188 2580 8192
rect 2516 8132 2520 8188
rect 2520 8132 2576 8188
rect 2576 8132 2580 8188
rect 2516 8128 2580 8132
rect 2596 8188 2660 8192
rect 2596 8132 2600 8188
rect 2600 8132 2656 8188
rect 2656 8132 2660 8188
rect 2596 8128 2660 8132
rect 2676 8188 2740 8192
rect 2676 8132 2680 8188
rect 2680 8132 2736 8188
rect 2736 8132 2740 8188
rect 2676 8128 2740 8132
rect 2756 8188 2820 8192
rect 2756 8132 2760 8188
rect 2760 8132 2816 8188
rect 2816 8132 2820 8188
rect 2756 8128 2820 8132
rect 5644 8188 5708 8192
rect 5644 8132 5648 8188
rect 5648 8132 5704 8188
rect 5704 8132 5708 8188
rect 5644 8128 5708 8132
rect 5724 8188 5788 8192
rect 5724 8132 5728 8188
rect 5728 8132 5784 8188
rect 5784 8132 5788 8188
rect 5724 8128 5788 8132
rect 5804 8188 5868 8192
rect 5804 8132 5808 8188
rect 5808 8132 5864 8188
rect 5864 8132 5868 8188
rect 5804 8128 5868 8132
rect 5884 8188 5948 8192
rect 5884 8132 5888 8188
rect 5888 8132 5944 8188
rect 5944 8132 5948 8188
rect 5884 8128 5948 8132
rect 8772 8188 8836 8192
rect 8772 8132 8776 8188
rect 8776 8132 8832 8188
rect 8832 8132 8836 8188
rect 8772 8128 8836 8132
rect 8852 8188 8916 8192
rect 8852 8132 8856 8188
rect 8856 8132 8912 8188
rect 8912 8132 8916 8188
rect 8852 8128 8916 8132
rect 8932 8188 8996 8192
rect 8932 8132 8936 8188
rect 8936 8132 8992 8188
rect 8992 8132 8996 8188
rect 8932 8128 8996 8132
rect 9012 8188 9076 8192
rect 9012 8132 9016 8188
rect 9016 8132 9072 8188
rect 9072 8132 9076 8188
rect 9012 8128 9076 8132
rect 11900 8188 11964 8192
rect 11900 8132 11904 8188
rect 11904 8132 11960 8188
rect 11960 8132 11964 8188
rect 11900 8128 11964 8132
rect 11980 8188 12044 8192
rect 11980 8132 11984 8188
rect 11984 8132 12040 8188
rect 12040 8132 12044 8188
rect 11980 8128 12044 8132
rect 12060 8188 12124 8192
rect 12060 8132 12064 8188
rect 12064 8132 12120 8188
rect 12120 8132 12124 8188
rect 12060 8128 12124 8132
rect 12140 8188 12204 8192
rect 12140 8132 12144 8188
rect 12144 8132 12200 8188
rect 12200 8132 12204 8188
rect 12140 8128 12204 8132
rect 4080 7644 4144 7648
rect 4080 7588 4084 7644
rect 4084 7588 4140 7644
rect 4140 7588 4144 7644
rect 4080 7584 4144 7588
rect 4160 7644 4224 7648
rect 4160 7588 4164 7644
rect 4164 7588 4220 7644
rect 4220 7588 4224 7644
rect 4160 7584 4224 7588
rect 4240 7644 4304 7648
rect 4240 7588 4244 7644
rect 4244 7588 4300 7644
rect 4300 7588 4304 7644
rect 4240 7584 4304 7588
rect 4320 7644 4384 7648
rect 4320 7588 4324 7644
rect 4324 7588 4380 7644
rect 4380 7588 4384 7644
rect 4320 7584 4384 7588
rect 7208 7644 7272 7648
rect 7208 7588 7212 7644
rect 7212 7588 7268 7644
rect 7268 7588 7272 7644
rect 7208 7584 7272 7588
rect 7288 7644 7352 7648
rect 7288 7588 7292 7644
rect 7292 7588 7348 7644
rect 7348 7588 7352 7644
rect 7288 7584 7352 7588
rect 7368 7644 7432 7648
rect 7368 7588 7372 7644
rect 7372 7588 7428 7644
rect 7428 7588 7432 7644
rect 7368 7584 7432 7588
rect 7448 7644 7512 7648
rect 7448 7588 7452 7644
rect 7452 7588 7508 7644
rect 7508 7588 7512 7644
rect 7448 7584 7512 7588
rect 10336 7644 10400 7648
rect 10336 7588 10340 7644
rect 10340 7588 10396 7644
rect 10396 7588 10400 7644
rect 10336 7584 10400 7588
rect 10416 7644 10480 7648
rect 10416 7588 10420 7644
rect 10420 7588 10476 7644
rect 10476 7588 10480 7644
rect 10416 7584 10480 7588
rect 10496 7644 10560 7648
rect 10496 7588 10500 7644
rect 10500 7588 10556 7644
rect 10556 7588 10560 7644
rect 10496 7584 10560 7588
rect 10576 7644 10640 7648
rect 10576 7588 10580 7644
rect 10580 7588 10636 7644
rect 10636 7588 10640 7644
rect 10576 7584 10640 7588
rect 2516 7100 2580 7104
rect 2516 7044 2520 7100
rect 2520 7044 2576 7100
rect 2576 7044 2580 7100
rect 2516 7040 2580 7044
rect 2596 7100 2660 7104
rect 2596 7044 2600 7100
rect 2600 7044 2656 7100
rect 2656 7044 2660 7100
rect 2596 7040 2660 7044
rect 2676 7100 2740 7104
rect 2676 7044 2680 7100
rect 2680 7044 2736 7100
rect 2736 7044 2740 7100
rect 2676 7040 2740 7044
rect 2756 7100 2820 7104
rect 2756 7044 2760 7100
rect 2760 7044 2816 7100
rect 2816 7044 2820 7100
rect 2756 7040 2820 7044
rect 5644 7100 5708 7104
rect 5644 7044 5648 7100
rect 5648 7044 5704 7100
rect 5704 7044 5708 7100
rect 5644 7040 5708 7044
rect 5724 7100 5788 7104
rect 5724 7044 5728 7100
rect 5728 7044 5784 7100
rect 5784 7044 5788 7100
rect 5724 7040 5788 7044
rect 5804 7100 5868 7104
rect 5804 7044 5808 7100
rect 5808 7044 5864 7100
rect 5864 7044 5868 7100
rect 5804 7040 5868 7044
rect 5884 7100 5948 7104
rect 5884 7044 5888 7100
rect 5888 7044 5944 7100
rect 5944 7044 5948 7100
rect 5884 7040 5948 7044
rect 8772 7100 8836 7104
rect 8772 7044 8776 7100
rect 8776 7044 8832 7100
rect 8832 7044 8836 7100
rect 8772 7040 8836 7044
rect 8852 7100 8916 7104
rect 8852 7044 8856 7100
rect 8856 7044 8912 7100
rect 8912 7044 8916 7100
rect 8852 7040 8916 7044
rect 8932 7100 8996 7104
rect 8932 7044 8936 7100
rect 8936 7044 8992 7100
rect 8992 7044 8996 7100
rect 8932 7040 8996 7044
rect 9012 7100 9076 7104
rect 9012 7044 9016 7100
rect 9016 7044 9072 7100
rect 9072 7044 9076 7100
rect 9012 7040 9076 7044
rect 11900 7100 11964 7104
rect 11900 7044 11904 7100
rect 11904 7044 11960 7100
rect 11960 7044 11964 7100
rect 11900 7040 11964 7044
rect 11980 7100 12044 7104
rect 11980 7044 11984 7100
rect 11984 7044 12040 7100
rect 12040 7044 12044 7100
rect 11980 7040 12044 7044
rect 12060 7100 12124 7104
rect 12060 7044 12064 7100
rect 12064 7044 12120 7100
rect 12120 7044 12124 7100
rect 12060 7040 12124 7044
rect 12140 7100 12204 7104
rect 12140 7044 12144 7100
rect 12144 7044 12200 7100
rect 12200 7044 12204 7100
rect 12140 7040 12204 7044
rect 4080 6556 4144 6560
rect 4080 6500 4084 6556
rect 4084 6500 4140 6556
rect 4140 6500 4144 6556
rect 4080 6496 4144 6500
rect 4160 6556 4224 6560
rect 4160 6500 4164 6556
rect 4164 6500 4220 6556
rect 4220 6500 4224 6556
rect 4160 6496 4224 6500
rect 4240 6556 4304 6560
rect 4240 6500 4244 6556
rect 4244 6500 4300 6556
rect 4300 6500 4304 6556
rect 4240 6496 4304 6500
rect 4320 6556 4384 6560
rect 4320 6500 4324 6556
rect 4324 6500 4380 6556
rect 4380 6500 4384 6556
rect 4320 6496 4384 6500
rect 7208 6556 7272 6560
rect 7208 6500 7212 6556
rect 7212 6500 7268 6556
rect 7268 6500 7272 6556
rect 7208 6496 7272 6500
rect 7288 6556 7352 6560
rect 7288 6500 7292 6556
rect 7292 6500 7348 6556
rect 7348 6500 7352 6556
rect 7288 6496 7352 6500
rect 7368 6556 7432 6560
rect 7368 6500 7372 6556
rect 7372 6500 7428 6556
rect 7428 6500 7432 6556
rect 7368 6496 7432 6500
rect 7448 6556 7512 6560
rect 7448 6500 7452 6556
rect 7452 6500 7508 6556
rect 7508 6500 7512 6556
rect 7448 6496 7512 6500
rect 10336 6556 10400 6560
rect 10336 6500 10340 6556
rect 10340 6500 10396 6556
rect 10396 6500 10400 6556
rect 10336 6496 10400 6500
rect 10416 6556 10480 6560
rect 10416 6500 10420 6556
rect 10420 6500 10476 6556
rect 10476 6500 10480 6556
rect 10416 6496 10480 6500
rect 10496 6556 10560 6560
rect 10496 6500 10500 6556
rect 10500 6500 10556 6556
rect 10556 6500 10560 6556
rect 10496 6496 10560 6500
rect 10576 6556 10640 6560
rect 10576 6500 10580 6556
rect 10580 6500 10636 6556
rect 10636 6500 10640 6556
rect 10576 6496 10640 6500
rect 2516 6012 2580 6016
rect 2516 5956 2520 6012
rect 2520 5956 2576 6012
rect 2576 5956 2580 6012
rect 2516 5952 2580 5956
rect 2596 6012 2660 6016
rect 2596 5956 2600 6012
rect 2600 5956 2656 6012
rect 2656 5956 2660 6012
rect 2596 5952 2660 5956
rect 2676 6012 2740 6016
rect 2676 5956 2680 6012
rect 2680 5956 2736 6012
rect 2736 5956 2740 6012
rect 2676 5952 2740 5956
rect 2756 6012 2820 6016
rect 2756 5956 2760 6012
rect 2760 5956 2816 6012
rect 2816 5956 2820 6012
rect 2756 5952 2820 5956
rect 5644 6012 5708 6016
rect 5644 5956 5648 6012
rect 5648 5956 5704 6012
rect 5704 5956 5708 6012
rect 5644 5952 5708 5956
rect 5724 6012 5788 6016
rect 5724 5956 5728 6012
rect 5728 5956 5784 6012
rect 5784 5956 5788 6012
rect 5724 5952 5788 5956
rect 5804 6012 5868 6016
rect 5804 5956 5808 6012
rect 5808 5956 5864 6012
rect 5864 5956 5868 6012
rect 5804 5952 5868 5956
rect 5884 6012 5948 6016
rect 5884 5956 5888 6012
rect 5888 5956 5944 6012
rect 5944 5956 5948 6012
rect 5884 5952 5948 5956
rect 8772 6012 8836 6016
rect 8772 5956 8776 6012
rect 8776 5956 8832 6012
rect 8832 5956 8836 6012
rect 8772 5952 8836 5956
rect 8852 6012 8916 6016
rect 8852 5956 8856 6012
rect 8856 5956 8912 6012
rect 8912 5956 8916 6012
rect 8852 5952 8916 5956
rect 8932 6012 8996 6016
rect 8932 5956 8936 6012
rect 8936 5956 8992 6012
rect 8992 5956 8996 6012
rect 8932 5952 8996 5956
rect 9012 6012 9076 6016
rect 9012 5956 9016 6012
rect 9016 5956 9072 6012
rect 9072 5956 9076 6012
rect 9012 5952 9076 5956
rect 11900 6012 11964 6016
rect 11900 5956 11904 6012
rect 11904 5956 11960 6012
rect 11960 5956 11964 6012
rect 11900 5952 11964 5956
rect 11980 6012 12044 6016
rect 11980 5956 11984 6012
rect 11984 5956 12040 6012
rect 12040 5956 12044 6012
rect 11980 5952 12044 5956
rect 12060 6012 12124 6016
rect 12060 5956 12064 6012
rect 12064 5956 12120 6012
rect 12120 5956 12124 6012
rect 12060 5952 12124 5956
rect 12140 6012 12204 6016
rect 12140 5956 12144 6012
rect 12144 5956 12200 6012
rect 12200 5956 12204 6012
rect 12140 5952 12204 5956
rect 4080 5468 4144 5472
rect 4080 5412 4084 5468
rect 4084 5412 4140 5468
rect 4140 5412 4144 5468
rect 4080 5408 4144 5412
rect 4160 5468 4224 5472
rect 4160 5412 4164 5468
rect 4164 5412 4220 5468
rect 4220 5412 4224 5468
rect 4160 5408 4224 5412
rect 4240 5468 4304 5472
rect 4240 5412 4244 5468
rect 4244 5412 4300 5468
rect 4300 5412 4304 5468
rect 4240 5408 4304 5412
rect 4320 5468 4384 5472
rect 4320 5412 4324 5468
rect 4324 5412 4380 5468
rect 4380 5412 4384 5468
rect 4320 5408 4384 5412
rect 7208 5468 7272 5472
rect 7208 5412 7212 5468
rect 7212 5412 7268 5468
rect 7268 5412 7272 5468
rect 7208 5408 7272 5412
rect 7288 5468 7352 5472
rect 7288 5412 7292 5468
rect 7292 5412 7348 5468
rect 7348 5412 7352 5468
rect 7288 5408 7352 5412
rect 7368 5468 7432 5472
rect 7368 5412 7372 5468
rect 7372 5412 7428 5468
rect 7428 5412 7432 5468
rect 7368 5408 7432 5412
rect 7448 5468 7512 5472
rect 7448 5412 7452 5468
rect 7452 5412 7508 5468
rect 7508 5412 7512 5468
rect 7448 5408 7512 5412
rect 10336 5468 10400 5472
rect 10336 5412 10340 5468
rect 10340 5412 10396 5468
rect 10396 5412 10400 5468
rect 10336 5408 10400 5412
rect 10416 5468 10480 5472
rect 10416 5412 10420 5468
rect 10420 5412 10476 5468
rect 10476 5412 10480 5468
rect 10416 5408 10480 5412
rect 10496 5468 10560 5472
rect 10496 5412 10500 5468
rect 10500 5412 10556 5468
rect 10556 5412 10560 5468
rect 10496 5408 10560 5412
rect 10576 5468 10640 5472
rect 10576 5412 10580 5468
rect 10580 5412 10636 5468
rect 10636 5412 10640 5468
rect 10576 5408 10640 5412
rect 2516 4924 2580 4928
rect 2516 4868 2520 4924
rect 2520 4868 2576 4924
rect 2576 4868 2580 4924
rect 2516 4864 2580 4868
rect 2596 4924 2660 4928
rect 2596 4868 2600 4924
rect 2600 4868 2656 4924
rect 2656 4868 2660 4924
rect 2596 4864 2660 4868
rect 2676 4924 2740 4928
rect 2676 4868 2680 4924
rect 2680 4868 2736 4924
rect 2736 4868 2740 4924
rect 2676 4864 2740 4868
rect 2756 4924 2820 4928
rect 2756 4868 2760 4924
rect 2760 4868 2816 4924
rect 2816 4868 2820 4924
rect 2756 4864 2820 4868
rect 5644 4924 5708 4928
rect 5644 4868 5648 4924
rect 5648 4868 5704 4924
rect 5704 4868 5708 4924
rect 5644 4864 5708 4868
rect 5724 4924 5788 4928
rect 5724 4868 5728 4924
rect 5728 4868 5784 4924
rect 5784 4868 5788 4924
rect 5724 4864 5788 4868
rect 5804 4924 5868 4928
rect 5804 4868 5808 4924
rect 5808 4868 5864 4924
rect 5864 4868 5868 4924
rect 5804 4864 5868 4868
rect 5884 4924 5948 4928
rect 5884 4868 5888 4924
rect 5888 4868 5944 4924
rect 5944 4868 5948 4924
rect 5884 4864 5948 4868
rect 8772 4924 8836 4928
rect 8772 4868 8776 4924
rect 8776 4868 8832 4924
rect 8832 4868 8836 4924
rect 8772 4864 8836 4868
rect 8852 4924 8916 4928
rect 8852 4868 8856 4924
rect 8856 4868 8912 4924
rect 8912 4868 8916 4924
rect 8852 4864 8916 4868
rect 8932 4924 8996 4928
rect 8932 4868 8936 4924
rect 8936 4868 8992 4924
rect 8992 4868 8996 4924
rect 8932 4864 8996 4868
rect 9012 4924 9076 4928
rect 9012 4868 9016 4924
rect 9016 4868 9072 4924
rect 9072 4868 9076 4924
rect 9012 4864 9076 4868
rect 11900 4924 11964 4928
rect 11900 4868 11904 4924
rect 11904 4868 11960 4924
rect 11960 4868 11964 4924
rect 11900 4864 11964 4868
rect 11980 4924 12044 4928
rect 11980 4868 11984 4924
rect 11984 4868 12040 4924
rect 12040 4868 12044 4924
rect 11980 4864 12044 4868
rect 12060 4924 12124 4928
rect 12060 4868 12064 4924
rect 12064 4868 12120 4924
rect 12120 4868 12124 4924
rect 12060 4864 12124 4868
rect 12140 4924 12204 4928
rect 12140 4868 12144 4924
rect 12144 4868 12200 4924
rect 12200 4868 12204 4924
rect 12140 4864 12204 4868
rect 4080 4380 4144 4384
rect 4080 4324 4084 4380
rect 4084 4324 4140 4380
rect 4140 4324 4144 4380
rect 4080 4320 4144 4324
rect 4160 4380 4224 4384
rect 4160 4324 4164 4380
rect 4164 4324 4220 4380
rect 4220 4324 4224 4380
rect 4160 4320 4224 4324
rect 4240 4380 4304 4384
rect 4240 4324 4244 4380
rect 4244 4324 4300 4380
rect 4300 4324 4304 4380
rect 4240 4320 4304 4324
rect 4320 4380 4384 4384
rect 4320 4324 4324 4380
rect 4324 4324 4380 4380
rect 4380 4324 4384 4380
rect 4320 4320 4384 4324
rect 7208 4380 7272 4384
rect 7208 4324 7212 4380
rect 7212 4324 7268 4380
rect 7268 4324 7272 4380
rect 7208 4320 7272 4324
rect 7288 4380 7352 4384
rect 7288 4324 7292 4380
rect 7292 4324 7348 4380
rect 7348 4324 7352 4380
rect 7288 4320 7352 4324
rect 7368 4380 7432 4384
rect 7368 4324 7372 4380
rect 7372 4324 7428 4380
rect 7428 4324 7432 4380
rect 7368 4320 7432 4324
rect 7448 4380 7512 4384
rect 7448 4324 7452 4380
rect 7452 4324 7508 4380
rect 7508 4324 7512 4380
rect 7448 4320 7512 4324
rect 10336 4380 10400 4384
rect 10336 4324 10340 4380
rect 10340 4324 10396 4380
rect 10396 4324 10400 4380
rect 10336 4320 10400 4324
rect 10416 4380 10480 4384
rect 10416 4324 10420 4380
rect 10420 4324 10476 4380
rect 10476 4324 10480 4380
rect 10416 4320 10480 4324
rect 10496 4380 10560 4384
rect 10496 4324 10500 4380
rect 10500 4324 10556 4380
rect 10556 4324 10560 4380
rect 10496 4320 10560 4324
rect 10576 4380 10640 4384
rect 10576 4324 10580 4380
rect 10580 4324 10636 4380
rect 10636 4324 10640 4380
rect 10576 4320 10640 4324
rect 2516 3836 2580 3840
rect 2516 3780 2520 3836
rect 2520 3780 2576 3836
rect 2576 3780 2580 3836
rect 2516 3776 2580 3780
rect 2596 3836 2660 3840
rect 2596 3780 2600 3836
rect 2600 3780 2656 3836
rect 2656 3780 2660 3836
rect 2596 3776 2660 3780
rect 2676 3836 2740 3840
rect 2676 3780 2680 3836
rect 2680 3780 2736 3836
rect 2736 3780 2740 3836
rect 2676 3776 2740 3780
rect 2756 3836 2820 3840
rect 2756 3780 2760 3836
rect 2760 3780 2816 3836
rect 2816 3780 2820 3836
rect 2756 3776 2820 3780
rect 5644 3836 5708 3840
rect 5644 3780 5648 3836
rect 5648 3780 5704 3836
rect 5704 3780 5708 3836
rect 5644 3776 5708 3780
rect 5724 3836 5788 3840
rect 5724 3780 5728 3836
rect 5728 3780 5784 3836
rect 5784 3780 5788 3836
rect 5724 3776 5788 3780
rect 5804 3836 5868 3840
rect 5804 3780 5808 3836
rect 5808 3780 5864 3836
rect 5864 3780 5868 3836
rect 5804 3776 5868 3780
rect 5884 3836 5948 3840
rect 5884 3780 5888 3836
rect 5888 3780 5944 3836
rect 5944 3780 5948 3836
rect 5884 3776 5948 3780
rect 8772 3836 8836 3840
rect 8772 3780 8776 3836
rect 8776 3780 8832 3836
rect 8832 3780 8836 3836
rect 8772 3776 8836 3780
rect 8852 3836 8916 3840
rect 8852 3780 8856 3836
rect 8856 3780 8912 3836
rect 8912 3780 8916 3836
rect 8852 3776 8916 3780
rect 8932 3836 8996 3840
rect 8932 3780 8936 3836
rect 8936 3780 8992 3836
rect 8992 3780 8996 3836
rect 8932 3776 8996 3780
rect 9012 3836 9076 3840
rect 9012 3780 9016 3836
rect 9016 3780 9072 3836
rect 9072 3780 9076 3836
rect 9012 3776 9076 3780
rect 11900 3836 11964 3840
rect 11900 3780 11904 3836
rect 11904 3780 11960 3836
rect 11960 3780 11964 3836
rect 11900 3776 11964 3780
rect 11980 3836 12044 3840
rect 11980 3780 11984 3836
rect 11984 3780 12040 3836
rect 12040 3780 12044 3836
rect 11980 3776 12044 3780
rect 12060 3836 12124 3840
rect 12060 3780 12064 3836
rect 12064 3780 12120 3836
rect 12120 3780 12124 3836
rect 12060 3776 12124 3780
rect 12140 3836 12204 3840
rect 12140 3780 12144 3836
rect 12144 3780 12200 3836
rect 12200 3780 12204 3836
rect 12140 3776 12204 3780
rect 4080 3292 4144 3296
rect 4080 3236 4084 3292
rect 4084 3236 4140 3292
rect 4140 3236 4144 3292
rect 4080 3232 4144 3236
rect 4160 3292 4224 3296
rect 4160 3236 4164 3292
rect 4164 3236 4220 3292
rect 4220 3236 4224 3292
rect 4160 3232 4224 3236
rect 4240 3292 4304 3296
rect 4240 3236 4244 3292
rect 4244 3236 4300 3292
rect 4300 3236 4304 3292
rect 4240 3232 4304 3236
rect 4320 3292 4384 3296
rect 4320 3236 4324 3292
rect 4324 3236 4380 3292
rect 4380 3236 4384 3292
rect 4320 3232 4384 3236
rect 7208 3292 7272 3296
rect 7208 3236 7212 3292
rect 7212 3236 7268 3292
rect 7268 3236 7272 3292
rect 7208 3232 7272 3236
rect 7288 3292 7352 3296
rect 7288 3236 7292 3292
rect 7292 3236 7348 3292
rect 7348 3236 7352 3292
rect 7288 3232 7352 3236
rect 7368 3292 7432 3296
rect 7368 3236 7372 3292
rect 7372 3236 7428 3292
rect 7428 3236 7432 3292
rect 7368 3232 7432 3236
rect 7448 3292 7512 3296
rect 7448 3236 7452 3292
rect 7452 3236 7508 3292
rect 7508 3236 7512 3292
rect 7448 3232 7512 3236
rect 10336 3292 10400 3296
rect 10336 3236 10340 3292
rect 10340 3236 10396 3292
rect 10396 3236 10400 3292
rect 10336 3232 10400 3236
rect 10416 3292 10480 3296
rect 10416 3236 10420 3292
rect 10420 3236 10476 3292
rect 10476 3236 10480 3292
rect 10416 3232 10480 3236
rect 10496 3292 10560 3296
rect 10496 3236 10500 3292
rect 10500 3236 10556 3292
rect 10556 3236 10560 3292
rect 10496 3232 10560 3236
rect 10576 3292 10640 3296
rect 10576 3236 10580 3292
rect 10580 3236 10636 3292
rect 10636 3236 10640 3292
rect 10576 3232 10640 3236
rect 2516 2748 2580 2752
rect 2516 2692 2520 2748
rect 2520 2692 2576 2748
rect 2576 2692 2580 2748
rect 2516 2688 2580 2692
rect 2596 2748 2660 2752
rect 2596 2692 2600 2748
rect 2600 2692 2656 2748
rect 2656 2692 2660 2748
rect 2596 2688 2660 2692
rect 2676 2748 2740 2752
rect 2676 2692 2680 2748
rect 2680 2692 2736 2748
rect 2736 2692 2740 2748
rect 2676 2688 2740 2692
rect 2756 2748 2820 2752
rect 2756 2692 2760 2748
rect 2760 2692 2816 2748
rect 2816 2692 2820 2748
rect 2756 2688 2820 2692
rect 5644 2748 5708 2752
rect 5644 2692 5648 2748
rect 5648 2692 5704 2748
rect 5704 2692 5708 2748
rect 5644 2688 5708 2692
rect 5724 2748 5788 2752
rect 5724 2692 5728 2748
rect 5728 2692 5784 2748
rect 5784 2692 5788 2748
rect 5724 2688 5788 2692
rect 5804 2748 5868 2752
rect 5804 2692 5808 2748
rect 5808 2692 5864 2748
rect 5864 2692 5868 2748
rect 5804 2688 5868 2692
rect 5884 2748 5948 2752
rect 5884 2692 5888 2748
rect 5888 2692 5944 2748
rect 5944 2692 5948 2748
rect 5884 2688 5948 2692
rect 8772 2748 8836 2752
rect 8772 2692 8776 2748
rect 8776 2692 8832 2748
rect 8832 2692 8836 2748
rect 8772 2688 8836 2692
rect 8852 2748 8916 2752
rect 8852 2692 8856 2748
rect 8856 2692 8912 2748
rect 8912 2692 8916 2748
rect 8852 2688 8916 2692
rect 8932 2748 8996 2752
rect 8932 2692 8936 2748
rect 8936 2692 8992 2748
rect 8992 2692 8996 2748
rect 8932 2688 8996 2692
rect 9012 2748 9076 2752
rect 9012 2692 9016 2748
rect 9016 2692 9072 2748
rect 9072 2692 9076 2748
rect 9012 2688 9076 2692
rect 11900 2748 11964 2752
rect 11900 2692 11904 2748
rect 11904 2692 11960 2748
rect 11960 2692 11964 2748
rect 11900 2688 11964 2692
rect 11980 2748 12044 2752
rect 11980 2692 11984 2748
rect 11984 2692 12040 2748
rect 12040 2692 12044 2748
rect 11980 2688 12044 2692
rect 12060 2748 12124 2752
rect 12060 2692 12064 2748
rect 12064 2692 12120 2748
rect 12120 2692 12124 2748
rect 12060 2688 12124 2692
rect 12140 2748 12204 2752
rect 12140 2692 12144 2748
rect 12144 2692 12200 2748
rect 12200 2692 12204 2748
rect 12140 2688 12204 2692
rect 4080 2204 4144 2208
rect 4080 2148 4084 2204
rect 4084 2148 4140 2204
rect 4140 2148 4144 2204
rect 4080 2144 4144 2148
rect 4160 2204 4224 2208
rect 4160 2148 4164 2204
rect 4164 2148 4220 2204
rect 4220 2148 4224 2204
rect 4160 2144 4224 2148
rect 4240 2204 4304 2208
rect 4240 2148 4244 2204
rect 4244 2148 4300 2204
rect 4300 2148 4304 2204
rect 4240 2144 4304 2148
rect 4320 2204 4384 2208
rect 4320 2148 4324 2204
rect 4324 2148 4380 2204
rect 4380 2148 4384 2204
rect 4320 2144 4384 2148
rect 7208 2204 7272 2208
rect 7208 2148 7212 2204
rect 7212 2148 7268 2204
rect 7268 2148 7272 2204
rect 7208 2144 7272 2148
rect 7288 2204 7352 2208
rect 7288 2148 7292 2204
rect 7292 2148 7348 2204
rect 7348 2148 7352 2204
rect 7288 2144 7352 2148
rect 7368 2204 7432 2208
rect 7368 2148 7372 2204
rect 7372 2148 7428 2204
rect 7428 2148 7432 2204
rect 7368 2144 7432 2148
rect 7448 2204 7512 2208
rect 7448 2148 7452 2204
rect 7452 2148 7508 2204
rect 7508 2148 7512 2204
rect 7448 2144 7512 2148
rect 10336 2204 10400 2208
rect 10336 2148 10340 2204
rect 10340 2148 10396 2204
rect 10396 2148 10400 2204
rect 10336 2144 10400 2148
rect 10416 2204 10480 2208
rect 10416 2148 10420 2204
rect 10420 2148 10476 2204
rect 10476 2148 10480 2204
rect 10416 2144 10480 2148
rect 10496 2204 10560 2208
rect 10496 2148 10500 2204
rect 10500 2148 10556 2204
rect 10556 2148 10560 2204
rect 10496 2144 10560 2148
rect 10576 2204 10640 2208
rect 10576 2148 10580 2204
rect 10580 2148 10636 2204
rect 10636 2148 10640 2204
rect 10576 2144 10640 2148
<< metal4 >>
rect 2508 14720 2828 14736
rect 2508 14656 2516 14720
rect 2580 14656 2596 14720
rect 2660 14656 2676 14720
rect 2740 14656 2756 14720
rect 2820 14656 2828 14720
rect 2508 13632 2828 14656
rect 2508 13568 2516 13632
rect 2580 13568 2596 13632
rect 2660 13568 2676 13632
rect 2740 13568 2756 13632
rect 2820 13568 2828 13632
rect 2508 13194 2828 13568
rect 2508 12958 2550 13194
rect 2786 12958 2828 13194
rect 2508 12544 2828 12958
rect 2508 12480 2516 12544
rect 2580 12480 2596 12544
rect 2660 12480 2676 12544
rect 2740 12480 2756 12544
rect 2820 12480 2828 12544
rect 2508 11456 2828 12480
rect 2508 11392 2516 11456
rect 2580 11392 2596 11456
rect 2660 11392 2676 11456
rect 2740 11392 2756 11456
rect 2820 11392 2828 11456
rect 2508 10368 2828 11392
rect 2508 10304 2516 10368
rect 2580 10304 2596 10368
rect 2660 10304 2676 10368
rect 2740 10304 2756 10368
rect 2820 10304 2828 10368
rect 2508 10066 2828 10304
rect 2508 9830 2550 10066
rect 2786 9830 2828 10066
rect 2508 9280 2828 9830
rect 2508 9216 2516 9280
rect 2580 9216 2596 9280
rect 2660 9216 2676 9280
rect 2740 9216 2756 9280
rect 2820 9216 2828 9280
rect 2508 8192 2828 9216
rect 2508 8128 2516 8192
rect 2580 8128 2596 8192
rect 2660 8128 2676 8192
rect 2740 8128 2756 8192
rect 2820 8128 2828 8192
rect 2508 7104 2828 8128
rect 2508 7040 2516 7104
rect 2580 7040 2596 7104
rect 2660 7040 2676 7104
rect 2740 7040 2756 7104
rect 2820 7040 2828 7104
rect 2508 6938 2828 7040
rect 2508 6702 2550 6938
rect 2786 6702 2828 6938
rect 2508 6016 2828 6702
rect 2508 5952 2516 6016
rect 2580 5952 2596 6016
rect 2660 5952 2676 6016
rect 2740 5952 2756 6016
rect 2820 5952 2828 6016
rect 2508 4928 2828 5952
rect 2508 4864 2516 4928
rect 2580 4864 2596 4928
rect 2660 4864 2676 4928
rect 2740 4864 2756 4928
rect 2820 4864 2828 4928
rect 2508 3840 2828 4864
rect 2508 3776 2516 3840
rect 2580 3810 2596 3840
rect 2660 3810 2676 3840
rect 2740 3810 2756 3840
rect 2820 3776 2828 3840
rect 2508 3574 2550 3776
rect 2786 3574 2828 3776
rect 2508 2752 2828 3574
rect 2508 2688 2516 2752
rect 2580 2688 2596 2752
rect 2660 2688 2676 2752
rect 2740 2688 2756 2752
rect 2820 2688 2828 2752
rect 2508 2128 2828 2688
rect 4072 14176 4392 14736
rect 4072 14112 4080 14176
rect 4144 14112 4160 14176
rect 4224 14112 4240 14176
rect 4304 14112 4320 14176
rect 4384 14112 4392 14176
rect 4072 13088 4392 14112
rect 4072 13024 4080 13088
rect 4144 13024 4160 13088
rect 4224 13024 4240 13088
rect 4304 13024 4320 13088
rect 4384 13024 4392 13088
rect 4072 12000 4392 13024
rect 4072 11936 4080 12000
rect 4144 11936 4160 12000
rect 4224 11936 4240 12000
rect 4304 11936 4320 12000
rect 4384 11936 4392 12000
rect 4072 11630 4392 11936
rect 4072 11394 4114 11630
rect 4350 11394 4392 11630
rect 4072 10912 4392 11394
rect 4072 10848 4080 10912
rect 4144 10848 4160 10912
rect 4224 10848 4240 10912
rect 4304 10848 4320 10912
rect 4384 10848 4392 10912
rect 4072 9824 4392 10848
rect 4072 9760 4080 9824
rect 4144 9760 4160 9824
rect 4224 9760 4240 9824
rect 4304 9760 4320 9824
rect 4384 9760 4392 9824
rect 4072 8736 4392 9760
rect 4072 8672 4080 8736
rect 4144 8672 4160 8736
rect 4224 8672 4240 8736
rect 4304 8672 4320 8736
rect 4384 8672 4392 8736
rect 4072 8502 4392 8672
rect 4072 8266 4114 8502
rect 4350 8266 4392 8502
rect 4072 7648 4392 8266
rect 4072 7584 4080 7648
rect 4144 7584 4160 7648
rect 4224 7584 4240 7648
rect 4304 7584 4320 7648
rect 4384 7584 4392 7648
rect 4072 6560 4392 7584
rect 4072 6496 4080 6560
rect 4144 6496 4160 6560
rect 4224 6496 4240 6560
rect 4304 6496 4320 6560
rect 4384 6496 4392 6560
rect 4072 5472 4392 6496
rect 4072 5408 4080 5472
rect 4144 5408 4160 5472
rect 4224 5408 4240 5472
rect 4304 5408 4320 5472
rect 4384 5408 4392 5472
rect 4072 5374 4392 5408
rect 4072 5138 4114 5374
rect 4350 5138 4392 5374
rect 4072 4384 4392 5138
rect 4072 4320 4080 4384
rect 4144 4320 4160 4384
rect 4224 4320 4240 4384
rect 4304 4320 4320 4384
rect 4384 4320 4392 4384
rect 4072 3296 4392 4320
rect 4072 3232 4080 3296
rect 4144 3232 4160 3296
rect 4224 3232 4240 3296
rect 4304 3232 4320 3296
rect 4384 3232 4392 3296
rect 4072 2208 4392 3232
rect 4072 2144 4080 2208
rect 4144 2144 4160 2208
rect 4224 2144 4240 2208
rect 4304 2144 4320 2208
rect 4384 2144 4392 2208
rect 4072 2128 4392 2144
rect 5636 14720 5956 14736
rect 5636 14656 5644 14720
rect 5708 14656 5724 14720
rect 5788 14656 5804 14720
rect 5868 14656 5884 14720
rect 5948 14656 5956 14720
rect 5636 13632 5956 14656
rect 5636 13568 5644 13632
rect 5708 13568 5724 13632
rect 5788 13568 5804 13632
rect 5868 13568 5884 13632
rect 5948 13568 5956 13632
rect 5636 13194 5956 13568
rect 5636 12958 5678 13194
rect 5914 12958 5956 13194
rect 5636 12544 5956 12958
rect 5636 12480 5644 12544
rect 5708 12480 5724 12544
rect 5788 12480 5804 12544
rect 5868 12480 5884 12544
rect 5948 12480 5956 12544
rect 5636 11456 5956 12480
rect 5636 11392 5644 11456
rect 5708 11392 5724 11456
rect 5788 11392 5804 11456
rect 5868 11392 5884 11456
rect 5948 11392 5956 11456
rect 5636 10368 5956 11392
rect 5636 10304 5644 10368
rect 5708 10304 5724 10368
rect 5788 10304 5804 10368
rect 5868 10304 5884 10368
rect 5948 10304 5956 10368
rect 5636 10066 5956 10304
rect 5636 9830 5678 10066
rect 5914 9830 5956 10066
rect 5636 9280 5956 9830
rect 5636 9216 5644 9280
rect 5708 9216 5724 9280
rect 5788 9216 5804 9280
rect 5868 9216 5884 9280
rect 5948 9216 5956 9280
rect 5636 8192 5956 9216
rect 5636 8128 5644 8192
rect 5708 8128 5724 8192
rect 5788 8128 5804 8192
rect 5868 8128 5884 8192
rect 5948 8128 5956 8192
rect 5636 7104 5956 8128
rect 5636 7040 5644 7104
rect 5708 7040 5724 7104
rect 5788 7040 5804 7104
rect 5868 7040 5884 7104
rect 5948 7040 5956 7104
rect 5636 6938 5956 7040
rect 5636 6702 5678 6938
rect 5914 6702 5956 6938
rect 5636 6016 5956 6702
rect 5636 5952 5644 6016
rect 5708 5952 5724 6016
rect 5788 5952 5804 6016
rect 5868 5952 5884 6016
rect 5948 5952 5956 6016
rect 5636 4928 5956 5952
rect 5636 4864 5644 4928
rect 5708 4864 5724 4928
rect 5788 4864 5804 4928
rect 5868 4864 5884 4928
rect 5948 4864 5956 4928
rect 5636 3840 5956 4864
rect 5636 3776 5644 3840
rect 5708 3810 5724 3840
rect 5788 3810 5804 3840
rect 5868 3810 5884 3840
rect 5948 3776 5956 3840
rect 5636 3574 5678 3776
rect 5914 3574 5956 3776
rect 5636 2752 5956 3574
rect 5636 2688 5644 2752
rect 5708 2688 5724 2752
rect 5788 2688 5804 2752
rect 5868 2688 5884 2752
rect 5948 2688 5956 2752
rect 5636 2128 5956 2688
rect 7200 14176 7520 14736
rect 7200 14112 7208 14176
rect 7272 14112 7288 14176
rect 7352 14112 7368 14176
rect 7432 14112 7448 14176
rect 7512 14112 7520 14176
rect 7200 13088 7520 14112
rect 7200 13024 7208 13088
rect 7272 13024 7288 13088
rect 7352 13024 7368 13088
rect 7432 13024 7448 13088
rect 7512 13024 7520 13088
rect 7200 12000 7520 13024
rect 7200 11936 7208 12000
rect 7272 11936 7288 12000
rect 7352 11936 7368 12000
rect 7432 11936 7448 12000
rect 7512 11936 7520 12000
rect 7200 11630 7520 11936
rect 7200 11394 7242 11630
rect 7478 11394 7520 11630
rect 7200 10912 7520 11394
rect 7200 10848 7208 10912
rect 7272 10848 7288 10912
rect 7352 10848 7368 10912
rect 7432 10848 7448 10912
rect 7512 10848 7520 10912
rect 7200 9824 7520 10848
rect 7200 9760 7208 9824
rect 7272 9760 7288 9824
rect 7352 9760 7368 9824
rect 7432 9760 7448 9824
rect 7512 9760 7520 9824
rect 7200 8736 7520 9760
rect 7200 8672 7208 8736
rect 7272 8672 7288 8736
rect 7352 8672 7368 8736
rect 7432 8672 7448 8736
rect 7512 8672 7520 8736
rect 7200 8502 7520 8672
rect 7200 8266 7242 8502
rect 7478 8266 7520 8502
rect 7200 7648 7520 8266
rect 7200 7584 7208 7648
rect 7272 7584 7288 7648
rect 7352 7584 7368 7648
rect 7432 7584 7448 7648
rect 7512 7584 7520 7648
rect 7200 6560 7520 7584
rect 7200 6496 7208 6560
rect 7272 6496 7288 6560
rect 7352 6496 7368 6560
rect 7432 6496 7448 6560
rect 7512 6496 7520 6560
rect 7200 5472 7520 6496
rect 7200 5408 7208 5472
rect 7272 5408 7288 5472
rect 7352 5408 7368 5472
rect 7432 5408 7448 5472
rect 7512 5408 7520 5472
rect 7200 5374 7520 5408
rect 7200 5138 7242 5374
rect 7478 5138 7520 5374
rect 7200 4384 7520 5138
rect 7200 4320 7208 4384
rect 7272 4320 7288 4384
rect 7352 4320 7368 4384
rect 7432 4320 7448 4384
rect 7512 4320 7520 4384
rect 7200 3296 7520 4320
rect 7200 3232 7208 3296
rect 7272 3232 7288 3296
rect 7352 3232 7368 3296
rect 7432 3232 7448 3296
rect 7512 3232 7520 3296
rect 7200 2208 7520 3232
rect 7200 2144 7208 2208
rect 7272 2144 7288 2208
rect 7352 2144 7368 2208
rect 7432 2144 7448 2208
rect 7512 2144 7520 2208
rect 7200 2128 7520 2144
rect 8764 14720 9084 14736
rect 8764 14656 8772 14720
rect 8836 14656 8852 14720
rect 8916 14656 8932 14720
rect 8996 14656 9012 14720
rect 9076 14656 9084 14720
rect 8764 13632 9084 14656
rect 8764 13568 8772 13632
rect 8836 13568 8852 13632
rect 8916 13568 8932 13632
rect 8996 13568 9012 13632
rect 9076 13568 9084 13632
rect 8764 13194 9084 13568
rect 8764 12958 8806 13194
rect 9042 12958 9084 13194
rect 8764 12544 9084 12958
rect 8764 12480 8772 12544
rect 8836 12480 8852 12544
rect 8916 12480 8932 12544
rect 8996 12480 9012 12544
rect 9076 12480 9084 12544
rect 8764 11456 9084 12480
rect 8764 11392 8772 11456
rect 8836 11392 8852 11456
rect 8916 11392 8932 11456
rect 8996 11392 9012 11456
rect 9076 11392 9084 11456
rect 8764 10368 9084 11392
rect 8764 10304 8772 10368
rect 8836 10304 8852 10368
rect 8916 10304 8932 10368
rect 8996 10304 9012 10368
rect 9076 10304 9084 10368
rect 8764 10066 9084 10304
rect 8764 9830 8806 10066
rect 9042 9830 9084 10066
rect 8764 9280 9084 9830
rect 8764 9216 8772 9280
rect 8836 9216 8852 9280
rect 8916 9216 8932 9280
rect 8996 9216 9012 9280
rect 9076 9216 9084 9280
rect 8764 8192 9084 9216
rect 8764 8128 8772 8192
rect 8836 8128 8852 8192
rect 8916 8128 8932 8192
rect 8996 8128 9012 8192
rect 9076 8128 9084 8192
rect 8764 7104 9084 8128
rect 8764 7040 8772 7104
rect 8836 7040 8852 7104
rect 8916 7040 8932 7104
rect 8996 7040 9012 7104
rect 9076 7040 9084 7104
rect 8764 6938 9084 7040
rect 8764 6702 8806 6938
rect 9042 6702 9084 6938
rect 8764 6016 9084 6702
rect 8764 5952 8772 6016
rect 8836 5952 8852 6016
rect 8916 5952 8932 6016
rect 8996 5952 9012 6016
rect 9076 5952 9084 6016
rect 8764 4928 9084 5952
rect 8764 4864 8772 4928
rect 8836 4864 8852 4928
rect 8916 4864 8932 4928
rect 8996 4864 9012 4928
rect 9076 4864 9084 4928
rect 8764 3840 9084 4864
rect 8764 3776 8772 3840
rect 8836 3810 8852 3840
rect 8916 3810 8932 3840
rect 8996 3810 9012 3840
rect 9076 3776 9084 3840
rect 8764 3574 8806 3776
rect 9042 3574 9084 3776
rect 8764 2752 9084 3574
rect 8764 2688 8772 2752
rect 8836 2688 8852 2752
rect 8916 2688 8932 2752
rect 8996 2688 9012 2752
rect 9076 2688 9084 2752
rect 8764 2128 9084 2688
rect 10328 14176 10648 14736
rect 10328 14112 10336 14176
rect 10400 14112 10416 14176
rect 10480 14112 10496 14176
rect 10560 14112 10576 14176
rect 10640 14112 10648 14176
rect 10328 13088 10648 14112
rect 10328 13024 10336 13088
rect 10400 13024 10416 13088
rect 10480 13024 10496 13088
rect 10560 13024 10576 13088
rect 10640 13024 10648 13088
rect 10328 12000 10648 13024
rect 10328 11936 10336 12000
rect 10400 11936 10416 12000
rect 10480 11936 10496 12000
rect 10560 11936 10576 12000
rect 10640 11936 10648 12000
rect 10328 11630 10648 11936
rect 10328 11394 10370 11630
rect 10606 11394 10648 11630
rect 10328 10912 10648 11394
rect 10328 10848 10336 10912
rect 10400 10848 10416 10912
rect 10480 10848 10496 10912
rect 10560 10848 10576 10912
rect 10640 10848 10648 10912
rect 10328 9824 10648 10848
rect 10328 9760 10336 9824
rect 10400 9760 10416 9824
rect 10480 9760 10496 9824
rect 10560 9760 10576 9824
rect 10640 9760 10648 9824
rect 10328 8736 10648 9760
rect 10328 8672 10336 8736
rect 10400 8672 10416 8736
rect 10480 8672 10496 8736
rect 10560 8672 10576 8736
rect 10640 8672 10648 8736
rect 10328 8502 10648 8672
rect 10328 8266 10370 8502
rect 10606 8266 10648 8502
rect 10328 7648 10648 8266
rect 10328 7584 10336 7648
rect 10400 7584 10416 7648
rect 10480 7584 10496 7648
rect 10560 7584 10576 7648
rect 10640 7584 10648 7648
rect 10328 6560 10648 7584
rect 10328 6496 10336 6560
rect 10400 6496 10416 6560
rect 10480 6496 10496 6560
rect 10560 6496 10576 6560
rect 10640 6496 10648 6560
rect 10328 5472 10648 6496
rect 10328 5408 10336 5472
rect 10400 5408 10416 5472
rect 10480 5408 10496 5472
rect 10560 5408 10576 5472
rect 10640 5408 10648 5472
rect 10328 5374 10648 5408
rect 10328 5138 10370 5374
rect 10606 5138 10648 5374
rect 10328 4384 10648 5138
rect 10328 4320 10336 4384
rect 10400 4320 10416 4384
rect 10480 4320 10496 4384
rect 10560 4320 10576 4384
rect 10640 4320 10648 4384
rect 10328 3296 10648 4320
rect 10328 3232 10336 3296
rect 10400 3232 10416 3296
rect 10480 3232 10496 3296
rect 10560 3232 10576 3296
rect 10640 3232 10648 3296
rect 10328 2208 10648 3232
rect 10328 2144 10336 2208
rect 10400 2144 10416 2208
rect 10480 2144 10496 2208
rect 10560 2144 10576 2208
rect 10640 2144 10648 2208
rect 10328 2128 10648 2144
rect 11892 14720 12212 14736
rect 11892 14656 11900 14720
rect 11964 14656 11980 14720
rect 12044 14656 12060 14720
rect 12124 14656 12140 14720
rect 12204 14656 12212 14720
rect 11892 13632 12212 14656
rect 11892 13568 11900 13632
rect 11964 13568 11980 13632
rect 12044 13568 12060 13632
rect 12124 13568 12140 13632
rect 12204 13568 12212 13632
rect 11892 13194 12212 13568
rect 11892 12958 11934 13194
rect 12170 12958 12212 13194
rect 11892 12544 12212 12958
rect 11892 12480 11900 12544
rect 11964 12480 11980 12544
rect 12044 12480 12060 12544
rect 12124 12480 12140 12544
rect 12204 12480 12212 12544
rect 11892 11456 12212 12480
rect 11892 11392 11900 11456
rect 11964 11392 11980 11456
rect 12044 11392 12060 11456
rect 12124 11392 12140 11456
rect 12204 11392 12212 11456
rect 11892 10368 12212 11392
rect 11892 10304 11900 10368
rect 11964 10304 11980 10368
rect 12044 10304 12060 10368
rect 12124 10304 12140 10368
rect 12204 10304 12212 10368
rect 11892 10066 12212 10304
rect 11892 9830 11934 10066
rect 12170 9830 12212 10066
rect 11892 9280 12212 9830
rect 11892 9216 11900 9280
rect 11964 9216 11980 9280
rect 12044 9216 12060 9280
rect 12124 9216 12140 9280
rect 12204 9216 12212 9280
rect 11892 8192 12212 9216
rect 11892 8128 11900 8192
rect 11964 8128 11980 8192
rect 12044 8128 12060 8192
rect 12124 8128 12140 8192
rect 12204 8128 12212 8192
rect 11892 7104 12212 8128
rect 11892 7040 11900 7104
rect 11964 7040 11980 7104
rect 12044 7040 12060 7104
rect 12124 7040 12140 7104
rect 12204 7040 12212 7104
rect 11892 6938 12212 7040
rect 11892 6702 11934 6938
rect 12170 6702 12212 6938
rect 11892 6016 12212 6702
rect 11892 5952 11900 6016
rect 11964 5952 11980 6016
rect 12044 5952 12060 6016
rect 12124 5952 12140 6016
rect 12204 5952 12212 6016
rect 11892 4928 12212 5952
rect 11892 4864 11900 4928
rect 11964 4864 11980 4928
rect 12044 4864 12060 4928
rect 12124 4864 12140 4928
rect 12204 4864 12212 4928
rect 11892 3840 12212 4864
rect 11892 3776 11900 3840
rect 11964 3810 11980 3840
rect 12044 3810 12060 3840
rect 12124 3810 12140 3840
rect 12204 3776 12212 3840
rect 11892 3574 11934 3776
rect 12170 3574 12212 3776
rect 11892 2752 12212 3574
rect 11892 2688 11900 2752
rect 11964 2688 11980 2752
rect 12044 2688 12060 2752
rect 12124 2688 12140 2752
rect 12204 2688 12212 2752
rect 11892 2128 12212 2688
<< via4 >>
rect 2550 12958 2786 13194
rect 2550 9830 2786 10066
rect 2550 6702 2786 6938
rect 2550 3776 2580 3810
rect 2580 3776 2596 3810
rect 2596 3776 2660 3810
rect 2660 3776 2676 3810
rect 2676 3776 2740 3810
rect 2740 3776 2756 3810
rect 2756 3776 2786 3810
rect 2550 3574 2786 3776
rect 4114 11394 4350 11630
rect 4114 8266 4350 8502
rect 4114 5138 4350 5374
rect 5678 12958 5914 13194
rect 5678 9830 5914 10066
rect 5678 6702 5914 6938
rect 5678 3776 5708 3810
rect 5708 3776 5724 3810
rect 5724 3776 5788 3810
rect 5788 3776 5804 3810
rect 5804 3776 5868 3810
rect 5868 3776 5884 3810
rect 5884 3776 5914 3810
rect 5678 3574 5914 3776
rect 7242 11394 7478 11630
rect 7242 8266 7478 8502
rect 7242 5138 7478 5374
rect 8806 12958 9042 13194
rect 8806 9830 9042 10066
rect 8806 6702 9042 6938
rect 8806 3776 8836 3810
rect 8836 3776 8852 3810
rect 8852 3776 8916 3810
rect 8916 3776 8932 3810
rect 8932 3776 8996 3810
rect 8996 3776 9012 3810
rect 9012 3776 9042 3810
rect 8806 3574 9042 3776
rect 10370 11394 10606 11630
rect 10370 8266 10606 8502
rect 10370 5138 10606 5374
rect 11934 12958 12170 13194
rect 11934 9830 12170 10066
rect 11934 6702 12170 6938
rect 11934 3776 11964 3810
rect 11964 3776 11980 3810
rect 11980 3776 12044 3810
rect 12044 3776 12060 3810
rect 12060 3776 12124 3810
rect 12124 3776 12140 3810
rect 12140 3776 12170 3810
rect 11934 3574 12170 3776
<< metal5 >>
rect 1104 13194 13616 13236
rect 1104 12958 2550 13194
rect 2786 12958 5678 13194
rect 5914 12958 8806 13194
rect 9042 12958 11934 13194
rect 12170 12958 13616 13194
rect 1104 12916 13616 12958
rect 1104 11630 13616 11672
rect 1104 11394 4114 11630
rect 4350 11394 7242 11630
rect 7478 11394 10370 11630
rect 10606 11394 13616 11630
rect 1104 11352 13616 11394
rect 1104 10066 13616 10108
rect 1104 9830 2550 10066
rect 2786 9830 5678 10066
rect 5914 9830 8806 10066
rect 9042 9830 11934 10066
rect 12170 9830 13616 10066
rect 1104 9788 13616 9830
rect 1104 8502 13616 8544
rect 1104 8266 4114 8502
rect 4350 8266 7242 8502
rect 7478 8266 10370 8502
rect 10606 8266 13616 8502
rect 1104 8224 13616 8266
rect 1104 6938 13616 6980
rect 1104 6702 2550 6938
rect 2786 6702 5678 6938
rect 5914 6702 8806 6938
rect 9042 6702 11934 6938
rect 12170 6702 13616 6938
rect 1104 6660 13616 6702
rect 1104 5374 13616 5416
rect 1104 5138 4114 5374
rect 4350 5138 7242 5374
rect 7478 5138 10370 5374
rect 10606 5138 13616 5374
rect 1104 5096 13616 5138
rect 1104 3810 13616 3852
rect 1104 3574 2550 3810
rect 2786 3574 5678 3810
rect 5914 3574 8806 3810
rect 9042 3574 11934 3810
rect 12170 3574 13616 3810
rect 1104 3532 13616 3574
use sky130_fd_sc_hd__decap_4  FILLER_0_3
timestamp 0
transform 1 0 1380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11
timestamp 0
transform 1 0 2116 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19
timestamp 0
transform 1 0 2852 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24
timestamp 0
transform 1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29
timestamp 0
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40
timestamp 0
transform 1 0 4784 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52
timestamp 0
transform 1 0 5888 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 0
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_69
timestamp 0
transform 1 0 7452 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77
timestamp 0
transform 1 0 8188 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83
timestamp 0
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 0
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 0
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 0
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113
timestamp 0
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_119
timestamp 0
transform 1 0 12052 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_129
timestamp 0
transform 1 0 12972 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_7
timestamp 0
transform 1 0 1748 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_13
timestamp 0
transform 1 0 2300 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_34
timestamp 0
transform 1 0 4232 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_46
timestamp 0
transform 1 0 5336 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp 0
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_60
timestamp 0
transform 1 0 6624 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_68
timestamp 0
transform 1 0 7360 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_80
timestamp 0
transform 1 0 8464 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_92
timestamp 0
transform 1 0 9568 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_104
timestamp 0
transform 1 0 10672 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 0
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_125
timestamp 0
transform 1 0 12604 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_23
timestamp 0
transform 1 0 3220 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 0
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_32
timestamp 0
transform 1 0 4048 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_44
timestamp 0
transform 1 0 5152 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_50
timestamp 0
transform 1 0 5704 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_71
timestamp 0
transform 1 0 7636 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_80
timestamp 0
transform 1 0 8464 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_105
timestamp 0
transform 1 0 10764 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_117
timestamp 0
transform 1 0 11868 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_129
timestamp 0
transform 1 0 12972 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3
timestamp 0
transform 1 0 1380 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_18
timestamp 0
transform 1 0 2760 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_22
timestamp 0
transform 1 0 3128 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_43
timestamp 0
transform 1 0 5060 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 0
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_57
timestamp 0
transform 1 0 6348 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_68
timestamp 0
transform 1 0 7360 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_84
timestamp 0
transform 1 0 8832 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_108
timestamp 0
transform 1 0 11040 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 0
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_125
timestamp 0
transform 1 0 12604 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_129
timestamp 0
transform 1 0 12972 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_3
timestamp 0
transform 1 0 1380 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_4_14
timestamp 0
transform 1 0 2392 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_26
timestamp 0
transform 1 0 3496 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_32
timestamp 0
transform 1 0 4048 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_38
timestamp 0
transform 1 0 4600 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_59
timestamp 0
transform 1 0 6532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_71
timestamp 0
transform 1 0 7636 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 0
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_105
timestamp 0
transform 1 0 10764 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_129
timestamp 0
transform 1 0 12972 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 0
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 0
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_27
timestamp 0
transform 1 0 3588 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_38
timestamp 0
transform 1 0 4600 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_50
timestamp 0
transform 1 0 5704 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_5_57
timestamp 0
transform 1 0 6348 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_65
timestamp 0
transform 1 0 7084 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_86
timestamp 0
transform 1 0 9016 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_98
timestamp 0
transform 1 0 10120 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_106
timestamp 0
transform 1 0 10856 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_5_113
timestamp 0
transform 1 0 11500 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_129
timestamp 0
transform 1 0 12972 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 0
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 0
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 0
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_29
timestamp 0
transform 1 0 3772 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_39
timestamp 0
transform 1 0 4692 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_51
timestamp 0
transform 1 0 5796 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_63
timestamp 0
transform 1 0 6900 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_75
timestamp 0
transform 1 0 8004 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 0
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_85
timestamp 0
transform 1 0 8924 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_91
timestamp 0
transform 1 0 9476 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_101
timestamp 0
transform 1 0 10396 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_105
timestamp 0
transform 1 0 10764 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_114
timestamp 0
transform 1 0 11592 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_122
timestamp 0
transform 1 0 12328 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_128
timestamp 0
transform 1 0 12880 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_132
timestamp 0
transform 1 0 13248 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 0
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_15
timestamp 0
transform 1 0 2484 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_21
timestamp 0
transform 1 0 3036 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_42
timestamp 0
transform 1 0 4968 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_54
timestamp 0
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_57
timestamp 0
transform 1 0 6348 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 0
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 0
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 0
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 0
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 0
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 0
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_125
timestamp 0
transform 1 0 12604 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_8_3
timestamp 0
transform 1 0 1380 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_11
timestamp 0
transform 1 0 2116 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_22
timestamp 0
transform 1 0 3128 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_8_29
timestamp 0
transform 1 0 3772 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_51
timestamp 0
transform 1 0 5796 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_72
timestamp 0
transform 1 0 7728 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_85
timestamp 0
transform 1 0 8924 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_98
timestamp 0
transform 1 0 10120 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_122
timestamp 0
transform 1 0 12328 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_130
timestamp 0
transform 1 0 13064 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_23
timestamp 0
transform 1 0 3220 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_30
timestamp 0
transform 1 0 3864 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_37
timestamp 0
transform 1 0 4508 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_49
timestamp 0
transform 1 0 5612 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 0
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_77
timestamp 0
transform 1 0 8188 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_84
timestamp 0
transform 1 0 8832 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_108
timestamp 0
transform 1 0 11040 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_113
timestamp 0
transform 1 0 11500 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_121
timestamp 0
transform 1 0 12236 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_129
timestamp 0
transform 1 0 12972 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_7
timestamp 0
transform 1 0 1748 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_14
timestamp 0
transform 1 0 2392 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_26
timestamp 0
transform 1 0 3496 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_32
timestamp 0
transform 1 0 4048 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_44
timestamp 0
transform 1 0 5152 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_56
timestamp 0
transform 1 0 6256 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_68
timestamp 0
transform 1 0 7360 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_80
timestamp 0
transform 1 0 8464 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_105
timestamp 0
transform 1 0 10764 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_129
timestamp 0
transform 1 0 12972 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 0
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 0
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_27
timestamp 0
transform 1 0 3588 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_34
timestamp 0
transform 1 0 4232 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_46
timestamp 0
transform 1 0 5336 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_54
timestamp 0
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 0
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 0
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_81
timestamp 0
transform 1 0 8556 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_89
timestamp 0
transform 1 0 9292 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 0
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 0
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 0
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 0
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_129
timestamp 0
transform 1 0 12972 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 0
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_15
timestamp 0
transform 1 0 2484 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_24
timestamp 0
transform 1 0 3312 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_38
timestamp 0
transform 1 0 4600 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_62
timestamp 0
transform 1 0 6808 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_74
timestamp 0
transform 1 0 7912 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_82
timestamp 0
transform 1 0 8648 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 0
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 0
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_129
timestamp 0
transform 1 0 12972 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_3
timestamp 0
transform 1 0 1380 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_24
timestamp 0
transform 1 0 3312 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_30
timestamp 0
transform 1 0 3864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 0
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 0
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_57
timestamp 0
transform 1 0 6348 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_65
timestamp 0
transform 1 0 7084 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_77
timestamp 0
transform 1 0 8188 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_83
timestamp 0
transform 1 0 8740 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 0
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 0
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 0
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_113
timestamp 0
transform 1 0 11500 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_117
timestamp 0
transform 1 0 11868 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_121
timestamp 0
transform 1 0 12236 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 0
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 0
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 0
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_29
timestamp 0
transform 1 0 3772 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_38
timestamp 0
transform 1 0 4600 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_45
timestamp 0
transform 1 0 5244 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_51
timestamp 0
transform 1 0 5796 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_72
timestamp 0
transform 1 0 7728 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_85
timestamp 0
transform 1 0 8924 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_14_111
timestamp 0
transform 1 0 11316 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_128
timestamp 0
transform 1 0 12880 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_132
timestamp 0
transform 1 0 13248 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_3
timestamp 0
transform 1 0 1380 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_9
timestamp 0
transform 1 0 1932 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_30
timestamp 0
transform 1 0 3864 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_42
timestamp 0
transform 1 0 4968 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_54
timestamp 0
transform 1 0 6072 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 0
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_69
timestamp 0
transform 1 0 7452 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_73
timestamp 0
transform 1 0 7820 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_78
timestamp 0
transform 1 0 8280 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_90
timestamp 0
transform 1 0 9384 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_102
timestamp 0
transform 1 0 10488 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_110
timestamp 0
transform 1 0 11224 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 0
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_125
timestamp 0
transform 1 0 12604 0 -1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 0
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 0
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 0
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_37
timestamp 0
transform 1 0 4508 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_49
timestamp 0
transform 1 0 5612 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_57
timestamp 0
transform 1 0 6348 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_80
timestamp 0
transform 1 0 8464 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_85
timestamp 0
transform 1 0 8924 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_93
timestamp 0
transform 1 0 9660 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_105
timestamp 0
transform 1 0 10764 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_128
timestamp 0
transform 1 0 12880 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_132
timestamp 0
transform 1 0 13248 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_7
timestamp 0
transform 1 0 1748 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_13
timestamp 0
transform 1 0 2300 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_34
timestamp 0
transform 1 0 4232 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_46
timestamp 0
transform 1 0 5336 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_54
timestamp 0
transform 1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_57
timestamp 0
transform 1 0 6348 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_17_66
timestamp 0
transform 1 0 7176 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_74
timestamp 0
transform 1 0 7912 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_95
timestamp 0
transform 1 0 9844 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_107
timestamp 0
transform 1 0 10948 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 0
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 0
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_125
timestamp 0
transform 1 0 12604 0 -1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 0
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 0
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 0
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_29
timestamp 0
transform 1 0 3772 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_37
timestamp 0
transform 1 0 4508 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_58
timestamp 0
transform 1 0 6440 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_70
timestamp 0
transform 1 0 7544 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_82
timestamp 0
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_85
timestamp 0
transform 1 0 8924 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_91
timestamp 0
transform 1 0 9476 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_112
timestamp 0
transform 1 0 11408 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_124
timestamp 0
transform 1 0 12512 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_132
timestamp 0
transform 1 0 13248 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 0
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 0
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 0
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_39
timestamp 0
transform 1 0 4692 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_47
timestamp 0
transform 1 0 5428 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 0
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_63
timestamp 0
transform 1 0 6900 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_75
timestamp 0
transform 1 0 8004 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_87
timestamp 0
transform 1 0 9108 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_19_102
timestamp 0
transform 1 0 10488 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_110
timestamp 0
transform 1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_113
timestamp 0
transform 1 0 11500 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_119
timestamp 0
transform 1 0 12052 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_124
timestamp 0
transform 1 0 12512 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_132
timestamp 0
transform 1 0 13248 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 0
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 0
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 0
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_29
timestamp 0
transform 1 0 3772 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_51
timestamp 0
transform 1 0 5796 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_79
timestamp 0
transform 1 0 8372 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 0
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_105
timestamp 0
transform 1 0 10764 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_117
timestamp 0
transform 1 0 11868 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_129
timestamp 0
transform 1 0 12972 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 0
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 0
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_27
timestamp 0
transform 1 0 3588 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_33
timestamp 0
transform 1 0 4140 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_37
timestamp 0
transform 1 0 4508 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_49
timestamp 0
transform 1 0 5612 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 0
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_60
timestamp 0
transform 1 0 6624 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_72
timestamp 0
transform 1 0 7728 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_84
timestamp 0
transform 1 0 8832 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_91
timestamp 0
transform 1 0 9476 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_21_101
timestamp 0
transform 1 0 10396 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_109
timestamp 0
transform 1 0 11132 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 0
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_125
timestamp 0
transform 1 0 12604 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_22_7
timestamp 0
transform 1 0 1748 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_15
timestamp 0
transform 1 0 2484 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_20
timestamp 0
transform 1 0 2944 0 1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 0
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 0
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_53
timestamp 0
transform 1 0 5980 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_57
timestamp 0
transform 1 0 6348 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_63
timestamp 0
transform 1 0 6900 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_75
timestamp 0
transform 1 0 8004 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 0
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 0
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_97
timestamp 0
transform 1 0 10028 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_105
timestamp 0
transform 1 0 10764 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_111
timestamp 0
transform 1 0 11316 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_113
timestamp 0
transform 1 0 11500 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_129
timestamp 0
transform 1 0 12972 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 0
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 0
transform -1 0 13616 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 0
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 0
transform -1 0 13616 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 0
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 0
transform -1 0 13616 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 0
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 0
transform -1 0 13616 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 0
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 0
transform -1 0 13616 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 0
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 0
transform -1 0 13616 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 0
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 0
transform -1 0 13616 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 0
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 0
transform -1 0 13616 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 0
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 0
transform -1 0 13616 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 0
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 0
transform -1 0 13616 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 0
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 0
transform -1 0 13616 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 0
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 0
transform -1 0 13616 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 0
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 0
transform -1 0 13616 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 0
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 0
transform -1 0 13616 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 0
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 0
transform -1 0 13616 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 0
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 0
transform -1 0 13616 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 0
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 0
transform -1 0 13616 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 0
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 0
transform -1 0 13616 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 0
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 0
transform -1 0 13616 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 0
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 0
transform -1 0 13616 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 0
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 0
transform -1 0 13616 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 0
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 0
transform -1 0 13616 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 0
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 0
transform -1 0 13616 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 0
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 0
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 0
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 0
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 0
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 0
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 0
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 0
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 0
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 0
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 0
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 0
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 0
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 0
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 0
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 0
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 0
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 0
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 0
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 0
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 0
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 0
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 0
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 0
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 0
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 0
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 0
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 0
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 0
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 0
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 0
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 0
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 0
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 0
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 0
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 0
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 0
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 0
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 0
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 0
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 0
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 0
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 0
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 0
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 0
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 0
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 0
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 0
transform 1 0 6256 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 0
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 0
transform 1 0 11408 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__a211o_1  _33_
timestamp 0
transform 1 0 4784 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _34_
timestamp 0
transform 1 0 6348 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _35_
timestamp 0
transform -1 0 6624 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _36_
timestamp 0
transform -1 0 8280 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _37_
timestamp 0
transform 1 0 3864 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _38_
timestamp 0
transform 1 0 9200 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _39_
timestamp 0
transform 1 0 3772 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__o21ba_1  _40_
timestamp 0
transform 1 0 2576 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _41_
timestamp 0
transform 1 0 4968 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _42_
timestamp 0
transform 1 0 3864 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__o21ba_1  _43_
timestamp 0
transform 1 0 3864 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _44_
timestamp 0
transform 1 0 7728 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _45_
timestamp 0
transform 1 0 6900 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__o21ba_1  _46_
timestamp 0
transform 1 0 6624 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _47_
timestamp 0
transform -1 0 9384 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _48_
timestamp 0
transform -1 0 9660 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__o21ba_1  _49_
timestamp 0
transform 1 0 9752 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _50_
timestamp 0
transform 1 0 3772 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _51_
timestamp 0
transform -1 0 10120 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _52_
timestamp 0
transform -1 0 10396 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__o21ba_1  _53_
timestamp 0
transform 1 0 10856 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _54_
timestamp 0
transform -1 0 8832 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _55_
timestamp 0
transform 1 0 9660 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _56_
timestamp 0
transform 1 0 9200 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _57_
timestamp 0
transform -1 0 2760 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _58_
timestamp 0
transform -1 0 2392 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _59_
timestamp 0
transform 1 0 2300 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _60_
timestamp 0
transform 1 0 2116 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _61_
timestamp 0
transform 1 0 12052 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _62_
timestamp 0
transform 1 0 11960 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _63_
timestamp 0
transform 1 0 6532 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _64_
timestamp 0
transform 1 0 6348 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _65__40
timestamp 0
transform -1 0 4508 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_1  _65_
timestamp 0
transform 1 0 3864 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _66_
timestamp 0
transform 1 0 5888 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _67_
timestamp 0
transform -1 0 11040 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _68_
timestamp 0
transform 1 0 9200 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _69_
timestamp 0
transform 1 0 11040 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _70_
timestamp 0
transform -1 0 4232 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _71_
timestamp 0
transform 1 0 6532 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _72_
timestamp 0
transform 1 0 6624 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _73_
timestamp 0
transform -1 0 6532 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _74_
timestamp 0
transform 1 0 10488 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _75_
timestamp 0
transform 1 0 4968 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _76_
timestamp 0
transform 1 0 4600 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _77_
timestamp 0
transform 1 0 8004 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _78_
timestamp 0
transform 1 0 8924 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _79_
timestamp 0
transform -1 0 12972 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _80_
timestamp 0
transform 1 0 2392 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _81_
timestamp 0
transform -1 0 4968 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _82_
timestamp 0
transform 1 0 8924 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _83_
timestamp 0
transform 1 0 9568 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _84_
timestamp 0
transform 1 0 3220 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _85_
timestamp 0
transform 1 0 7176 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _86_
timestamp 0
transform 1 0 3956 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _87_
timestamp 0
transform 1 0 1472 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _88_
timestamp 0
transform 1 0 3956 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _89_
timestamp 0
transform 1 0 6348 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _90_
timestamp 0
transform 1 0 9476 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _91_
timestamp 0
transform -1 0 3864 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _92_
timestamp 0
transform 1 0 11132 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _93_
timestamp 0
transform 1 0 8924 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _94_
timestamp 0
transform 1 0 8924 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _95_
timestamp 0
transform -1 0 3220 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _96_
timestamp 0
transform 1 0 1380 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _97_
timestamp 0
transform 1 0 11132 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _98_
timestamp 0
transform 1 0 5796 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_2  input1
timestamp 0
transform 1 0 1748 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  input2
timestamp 0
transform 1 0 3956 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 0
transform -1 0 2944 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 0
transform 1 0 12696 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output5
timestamp 0
transform 1 0 12604 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output6
timestamp 0
transform -1 0 1748 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output7
timestamp 0
transform 1 0 12604 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output8
timestamp 0
transform 1 0 12604 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output9
timestamp 0
transform -1 0 6900 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output10
timestamp 0
transform 1 0 11684 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output11
timestamp 0
transform -1 0 10764 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output12
timestamp 0
transform -1 0 1748 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output13
timestamp 0
transform -1 0 1748 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output14
timestamp 0
transform 1 0 12604 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output15
timestamp 0
transform 1 0 7820 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output16
timestamp 0
transform -1 0 1748 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater17
timestamp 0
transform -1 0 10396 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater18
timestamp 0
transform -1 0 7360 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater19
timestamp 0
transform -1 0 10856 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater20
timestamp 0
transform -1 0 7084 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  repeater21
timestamp 0
transform 1 0 8556 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  repeater22
timestamp 0
transform -1 0 7452 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater23
timestamp 0
transform -1 0 12236 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater24
timestamp 0
transform -1 0 9660 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater25
timestamp 0
transform -1 0 12512 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater26
timestamp 0
transform -1 0 12972 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater27
timestamp 0
transform 1 0 12512 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  repeater28
timestamp 0
transform -1 0 12972 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  repeater29
timestamp 0
transform -1 0 7176 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater30
timestamp 0
transform -1 0 5244 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater31
timestamp 0
transform -1 0 4232 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater32
timestamp 0
transform -1 0 9660 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater33
timestamp 0
transform -1 0 3864 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater34
timestamp 0
transform 1 0 4232 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater35
timestamp 0
transform -1 0 4048 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater36
timestamp 0
transform -1 0 4048 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater37
timestamp 0
transform -1 0 4048 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater38
timestamp 0
transform -1 0 8464 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater39
timestamp 0
transform -1 0 3312 0 1 2176
box -38 -48 314 592
<< labels >>
rlabel metal3 s 13944 8848 14744 8968 4 B[0]
port 1 nsew
rlabel metal3 s 0 15648 800 15768 4 B[1]
port 2 nsew
rlabel metal3 s 13944 12928 14744 13048 4 B[2]
port 3 nsew
rlabel metal3 s 13944 688 14744 808 4 B[3]
port 4 nsew
rlabel metal2 s 6458 16088 6514 16888 4 B[4]
port 5 nsew
rlabel metal2 s 18 0 74 800 4 CompOut
port 6 nsew
rlabel metal2 s 11610 0 11666 800 4 SH
port 7 nsew
rlabel metal5 s 1104 5096 13616 5416 4 VGND
port 8 nsew
rlabel metal5 s 1104 8224 13616 8544 4 VGND
port 8 nsew
rlabel metal5 s 1104 11352 13616 11672 4 VGND
port 8 nsew
rlabel metal4 s 4072 2128 4392 14736 4 VGND
port 8 nsew
rlabel metal4 s 7200 2128 7520 14736 4 VGND
port 8 nsew
rlabel metal4 s 10328 2128 10648 14736 4 VGND
port 8 nsew
rlabel metal5 s 1104 3532 13616 3852 4 VPWR
port 9 nsew
rlabel metal5 s 1104 6660 13616 6980 4 VPWR
port 9 nsew
rlabel metal5 s 1104 9788 13616 10108 4 VPWR
port 9 nsew
rlabel metal5 s 1104 12916 13616 13236 4 VPWR
port 9 nsew
rlabel metal4 s 2508 2128 2828 14736 4 VPWR
port 9 nsew
rlabel metal4 s 5636 2128 5956 14736 4 VPWR
port 9 nsew
rlabel metal4 s 8764 2128 9084 14736 4 VPWR
port 9 nsew
rlabel metal4 s 11892 2128 12212 14736 4 VPWR
port 9 nsew
rlabel metal2 s 3882 0 3938 800 4 clock
port 10 nsew
rlabel metal2 s 10322 16088 10378 16888 4 dataOut[0]
port 11 nsew
rlabel metal3 s 0 3408 800 3528 4 dataOut[1]
port 12 nsew
rlabel metal3 s 0 7488 800 7608 4 dataOut[2]
port 13 nsew
rlabel metal2 s 14186 16088 14242 16888 4 dataOut[3]
port 14 nsew
rlabel metal2 s 7746 0 7802 800 4 dataOut[4]
port 15 nsew
rlabel metal3 s 0 11568 800 11688 4 nEndCnv
port 16 nsew
rlabel metal2 s 2594 16088 2650 16888 4 nStartCnv
port 17 nsew
rlabel metal3 s 13944 4768 14744 4888 4 reset
port 18 nsew
<< properties >>
string FIXED_BBOX 0 0 14744 16888
<< end >>
