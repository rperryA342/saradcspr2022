* SPICE3 file created from caparry.ext - technology: sky130A

.option scale=10000u

X0 B0 vcommon sky130_fd_pr__cap_mim_m3_1 l=1000 w=1000
X1 B2 vcommon sky130_fd_pr__cap_mim_m3_1 l=1000 w=1000
X2 B2 vcommon sky130_fd_pr__cap_mim_m3_1 l=1000 w=1000
X3 B2 vcommon sky130_fd_pr__cap_mim_m3_1 l=1000 w=1000
X4 B2 vcommon sky130_fd_pr__cap_mim_m3_1 l=1000 w=1000
X5 B1 vcommon sky130_fd_pr__cap_mim_m3_1 l=1000 w=1000
X6 B1 vcommon sky130_fd_pr__cap_mim_m3_1 l=1000 w=1000
X7 B3 vcommon sky130_fd_pr__cap_mim_m3_1 l=1000 w=1000
X8 B3 vcommon sky130_fd_pr__cap_mim_m3_1 l=1000 w=1000
X9 B3 vcommon sky130_fd_pr__cap_mim_m3_1 l=1000 w=1000
X10 B3 vcommon sky130_fd_pr__cap_mim_m3_1 l=1000 w=1000
X11 B3 vcommon sky130_fd_pr__cap_mim_m3_1 l=1000 w=1000
X12 B3 vcommon sky130_fd_pr__cap_mim_m3_1 l=1000 w=1000
X13 B3 vcommon sky130_fd_pr__cap_mim_m3_1 l=1000 w=1000
X14 B3 vcommon sky130_fd_pr__cap_mim_m3_1 l=1000 w=1000
X15 B4 vcommon sky130_fd_pr__cap_mim_m3_1 l=1000 w=1000
X16 B4 vcommon sky130_fd_pr__cap_mim_m3_1 l=1000 w=1000
X17 B4 vcommon sky130_fd_pr__cap_mim_m3_1 l=1000 w=1000
X18 B4 vcommon sky130_fd_pr__cap_mim_m3_1 l=1000 w=1000
X19 B4 vcommon sky130_fd_pr__cap_mim_m3_1 l=1000 w=1000
X20 B4 vcommon sky130_fd_pr__cap_mim_m3_1 l=1000 w=1000
X21 B4 vcommon sky130_fd_pr__cap_mim_m3_1 l=1000 w=1000
X22 B4 vcommon sky130_fd_pr__cap_mim_m3_1 l=1000 w=1000
X23 B4 vcommon sky130_fd_pr__cap_mim_m3_1 l=1000 w=1000
X24 B4 vcommon sky130_fd_pr__cap_mim_m3_1 l=1000 w=1000
X25 B4 vcommon sky130_fd_pr__cap_mim_m3_1 l=1000 w=1000
X26 B4 vcommon sky130_fd_pr__cap_mim_m3_1 l=1000 w=1000
X27 B4 vcommon sky130_fd_pr__cap_mim_m3_1 l=1000 w=1000
X28 B4 vcommon sky130_fd_pr__cap_mim_m3_1 l=1000 w=1000
X29 B4 vcommon sky130_fd_pr__cap_mim_m3_1 l=1000 w=1000
X30 B4 vcommon sky130_fd_pr__cap_mim_m3_1 l=1000 w=1000
C0 vcommon B0 9.48fF
C1 vcommon B3 76.33fF
C2 B1 vcommon 18.96fF
C3 vcommon B2 38.16fF
C4 vcommon B4 152.90fF
C5 vcommon SUB 101.49fF **FLOATING
C6 B4 SUB 12.51fF **FLOATING
C7 B3 SUB 6.03fF **FLOATING
C8 B2 SUB 2.69fF **FLOATING
