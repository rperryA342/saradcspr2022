magic
tech sky130A
timestamp 1650135350
<< metal3 >>
rect 1060 1470 1070 1480
rect 5 -115 105 250
rect 2015 -115 2115 250
<< metal4 >>
rect 465 -180 565 0
rect 1550 -180 1650 100
rect 515 -1395 525 -1385
use mimcap2C  mimcap2C_1
timestamp 1649877975
transform 1 0 5 0 1 -1295
box 0 -100 2115 1380
use mimcap2C  mimcap2C_0
timestamp 1649877975
transform 1 0 0 0 1 100
box 0 -100 2115 1380
<< labels >>
rlabel metal3 1065 1480 1065 1480 1 common
rlabel metal4 520 -1395 520 -1395 5 top4C
<< end >>
