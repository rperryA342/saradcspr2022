** sch_path: /home/rperry/xschem_skywater/sar_adc_design/saradc2022/dacblock.sch


.param vONE=2
.param AGND=1
.param rt=5n
.param pw=250n
.param t0=100n
.param t0r=t0+rt
.param t1=t0r+pw
.param t1r=t1+rt
.param t2=t1r+pw
.param t2r=t2+rt
.param t3=t2r+pw
.param t3r=t3+rt
.param t4=t3r+pw
.param t4r=t4+rt
.param t5=t4r+pw
.param t5r=t5+rt
.param t6=t5r+pw
.param t6r=t6+rt
.param t7=t6r+pw
.param t7r=t7+rt
.param b2d=VONE
.param b1d=0
.param b0d=VONE
.param vadc=(b2d/4)+(b1d/8)+(b0d/16)+AGND



**.subckt dacblock Vin AGND VREF SH B0 B1 B2
*.ipin Vin
*.ipin AGND
*.ipin VREF
*.ipin SH
*.ipin B0
*.ipin B1
*.ipin B2
Vmax VDD GND 2
XC1 Vcommon c1v sky130_fd_pr__cap_mim_m3_1 W=10 L=10 MF=1 m=1
Vmax1 Vin GND {vadc}
Vmax3 AGND GND 1
V4 SH GND DC 0 pwl (0n 0 {t0} 0 {t0r} 2 {t1} 2 {t1r} 0)
XC5 CompOut GND sky130_fd_pr__cap_mim_m3_1 W=10 L=10 MF=1 m=1
Vmax4 VREF GND 2
XC2 Vcommon c2v sky130_fd_pr__cap_mim_m3_1 W=10 L=10 MF=1 m=1
V1 B1 GND DC 0 pwl (0n 0 {t0} 0 {t0r} 2 {t1} 2 {t1r} 0 {t4} 0 {t4r} 2 {t5} 2 {t5r} {b1d})
x3 Vcommon AGND CompOut skywater_comparator
V3 B0 GND dc 0 pwl (0n 0 {t0} 0 {t0r} 2 {t1} 2 {t1r} 0 {t6} 0 {t6r} 2 {t7} 2 {t7r} {b0d})
V5 B2 GND DC 0 pwl (0n 0 {t0} 0 {t0r} 2 {t1} 2 {t1r} 0 {t2} 0 {t2r} 2 {t3} 2 {t3r} {b2d})
XC6 Vcommon c4v sky130_fd_pr__cap_mim_m3_1 W=10 L=10 MF=4 m=4
XC7 Vcommon c3v sky130_fd_pr__cap_mim_m3_1 W=10 L=10 MF=2 m=2
x1 c4v SH Vin AGND VREF AGND B2 4x1analogmux
x2 c3v SH Vin AGND VREF AGND B1 4x1analogmux
x4 c2v SH Vin AGND VREF AGND B0 4x1analogmux
x5 c1v Vin AGND SH 2x1analogmux
x6 AGND SH net1 analog_switch
Vswitch net1 Vcommon 0
XC3 AGND GND sky130_fd_pr__cap_mim_m3_1 W=10 L=10 MF=1 m=1
**** begin user architecture code


.include opamp_sky130.sp

.tran 0.1 2000n
.control
run
**plot i(Vswitch)
write dacpassgate_testcircuit_v2.raw
plot v(SH) v(B0)+2 v(B1)+4 v(B2)+6
plot v(Vin)  v(vCommon)
**plot v(AGND)
plot v(c1v) v(c2v)+2 v(c3v)+4 v(c4v)+6
plot v(CompOut)
.endc



** opencircuitdesign pdks install
.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt


**** end user architecture code
**.ends

* expanding   symbol:  skywater_comparator.sym # of pins=3
** sym_path: /home/rperry/xschem_skywater/sar_adc_design/saradc2022/skywater_comparator.sym
** sch_path: /home/rperry/xschem_skywater/sar_adc_design/saradc2022/skywater_comparator.sch
.subckt skywater_comparator  Vmin Vpos Y
*.ipin Vpos
*.ipin Vmin
*.opin Y
x1 Y net1 VDD GND not W_N=1 L_N=0.15 W_P=2 L_P=0.15 m=10
x2 Vmin Vpos net1 VDD GND opamp_sky130
.ends


* expanding   symbol:  4x1analogmux.sym # of pins=7
** sym_path: /home/rperry/xschem_skywater/sar_adc_design/saradc2022/4x1analogmux.sym
** sch_path: /home/rperry/xschem_skywater/sar_adc_design/saradc2022/4x1analogmux.sch
.subckt 4x1analogmux  Vout S1 A3 A2 A1 A0 S0
*.ipin A3
*.ipin A2
*.ipin A1
*.ipin A0
*.ipin S1
*.ipin S0
*.opin Vout
x2 net2 A1 A0 S0 2x1analogmux
x3 Vout net1 net2 S1 2x1analogmux
x1 net1 A3 A2 S0 2x1analogmux
.ends


* expanding   symbol:  2x1analogmux.sym # of pins=4
** sym_path: /home/rperry/xschem_skywater/sar_adc_design/saradc2022/2x1analogmux.sym
** sch_path: /home/rperry/xschem_skywater/sar_adc_design/saradc2022/2x1analogmux.sch
.subckt 2x1analogmux  Vout A1 A0 S
*.ipin S
*.opin Vout
*.ipin A1
*.ipin A0
x1 net1 A1 Vout S dacpassgate
x2 S A0 Vout net1 dacpassgate
x3 net1 S VCC VSS not W_N=1 L_N=0.15 W_P=2 L_P=0.15 m=1
.ends


* expanding   symbol:  analog_switch.sym # of pins=3
** sym_path: /home/rperry/xschem_skywater/sar_adc_design/saradc2022/analog_switch.sym
** sch_path: /home/rperry/xschem_skywater/sar_adc_design/saradc2022/analog_switch.sch
.subckt analog_switch  Vin S Vout
*.ipin S
*.ipin Vin
*.opin Vout
x1 net1 Vin Vout S dacpassgate
x2 net1 S VCC VSS not W_N=1 L_N=0.15 W_P=2 L_P=0.15 m=1
.ends


* expanding   symbol:  not.sym # of pins=2
** sym_path: /home/rperry/xschem_skywater/sar_adc_design/saradc2022/not.sym
** sch_path: /home/rperry/xschem_skywater/sar_adc_design/saradc2022/not.sch
.subckt not  y a  VCCPIN  VSSPIN      W_N=1 L_N=0.15 W_P=2 L_P=0.15
*.opin y
*.ipin a
XM1 y a VSSPIN VSSPIN sky130_fd_pr__nfet_01v8 L=L_N W=W_N nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 y a VCCPIN VCCPIN sky130_fd_pr__pfet_01v8 L=L_P W=W_P nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  dacpassgate.sym # of pins=4
** sym_path: /home/rperry/xschem_skywater/sar_adc_design/saradc2022/dacpassgate.sym
** sch_path: /home/rperry/xschem_skywater/sar_adc_design/saradc2022/dacpassgate.sch
.subckt dacpassgate  GP A Z GN
*.iopin A
*.iopin Z
*.ipin GP
*.ipin GN
XM1 Z GN A GND sky130_fd_pr__nfet_01v8 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=10 m=10
XM2 Z GP A VDD sky130_fd_pr__pfet_01v8 L=0.5 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=10 m=10
.ends

.GLOBAL GND
.GLOBAL VDD
.end
