* SPICE3 file created from caparry.ext - technology: sky130A

*.option scale=10000u

.subckt caparray vcommon B50 B0 B1 B2 B3 B4 

X50 B50 vcommon sky130_fd_pr__cap_mim_m3_1 l=100u w=100u
X0  B0 vcommon sky130_fd_pr__cap_mim_m3_1 l=100u w=100u
X1  B2 vcommon sky130_fd_pr__cap_mim_m3_1 l=100u w=100u
X2  B2 vcommon sky130_fd_pr__cap_mim_m3_1 l=100u w=100u
X3  B2 vcommon sky130_fd_pr__cap_mim_m3_1 l=100u w=100u
X4  B2 vcommon sky130_fd_pr__cap_mim_m3_1 l=100u w=100u
X5  B1 vcommon sky130_fd_pr__cap_mim_m3_1 l=100u w=100u
X6  B1 vcommon sky130_fd_pr__cap_mim_m3_1 l=100u w=100u
X7  B3 vcommon sky130_fd_pr__cap_mim_m3_1 l=100u w=100u
X8  B3 vcommon sky130_fd_pr__cap_mim_m3_1 l=100u w=100u
X9  B3 vcommon sky130_fd_pr__cap_mim_m3_1 l=100u w=100u
X10 B3 vcommon sky130_fd_pr__cap_mim_m3_1 l=100u w=100u
X11 B3 vcommon sky130_fd_pr__cap_mim_m3_1 l=100u w=100u
X12 B3 vcommon sky130_fd_pr__cap_mim_m3_1 l=100u w=100u
X13 B3 vcommon sky130_fd_pr__cap_mim_m3_1 l=100u w=100u
X14 B3 vcommon sky130_fd_pr__cap_mim_m3_1 l=100u w=100u
X15 B4 vcommon sky130_fd_pr__cap_mim_m3_1 l=100u w=100u
X16 B4 vcommon sky130_fd_pr__cap_mim_m3_1 l=100u w=100u
X17 B4 vcommon sky130_fd_pr__cap_mim_m3_1 l=100u w=100u
X18 B4 vcommon sky130_fd_pr__cap_mim_m3_1 l=100u w=100u
X19 B4 vcommon sky130_fd_pr__cap_mim_m3_1 l=100u w=100u
X20 B4 vcommon sky130_fd_pr__cap_mim_m3_1 l=100u w=100u
X21 B4 vcommon sky130_fd_pr__cap_mim_m3_1 l=100u w=100u
X22 B4 vcommon sky130_fd_pr__cap_mim_m3_1 l=100u w=100u
X23 B4 vcommon sky130_fd_pr__cap_mim_m3_1 l=100u w=100u
X24 B4 vcommon sky130_fd_pr__cap_mim_m3_1 l=100u w=100u
X25 B4 vcommon sky130_fd_pr__cap_mim_m3_1 l=100u w=100u
X26 B4 vcommon sky130_fd_pr__cap_mim_m3_1 l=100u w=100u
X27 B4 vcommon sky130_fd_pr__cap_mim_m3_1 l=100u w=100u
X28 B4 vcommon sky130_fd_pr__cap_mim_m3_1 l=100u w=100u
X29 B4 vcommon sky130_fd_pr__cap_mim_m3_1 l=100u w=100u
X30 B4 vcommon sky130_fd_pr__cap_mim_m3_1 l=100u w=100u

.ends
