magic
tech sky130A
timestamp 1650405858
<< nwell >>
rect -107 629 1438 2771
<< nmos >>
rect 81 368 181 547
rect 482 368 582 547
rect -187 -617 -87 -149
rect 347 -757 447 155
rect 1643 -674 1743 2056
<< pmos >>
rect 77 691 177 1307
rect 506 691 606 1307
rect 936 810 1036 2645
<< ndiff >>
rect 1537 1975 1643 2056
rect 1538 1911 1643 1975
rect 1538 1871 1563 1911
rect 1604 1871 1643 1911
rect 1538 1822 1643 1871
rect 1538 1782 1563 1822
rect 1604 1782 1643 1822
rect -21 523 81 547
rect -21 483 1 523
rect 42 483 81 523
rect -21 434 81 483
rect -21 394 1 434
rect 42 394 81 434
rect -21 368 81 394
rect 181 523 291 547
rect 181 483 220 523
rect 261 483 291 523
rect 181 428 291 483
rect 181 388 216 428
rect 257 388 291 428
rect 181 368 291 388
rect 380 523 482 547
rect 380 483 402 523
rect 443 483 482 523
rect 380 434 482 483
rect 380 394 402 434
rect 443 394 482 434
rect 380 368 482 394
rect 582 523 692 547
rect 582 483 621 523
rect 662 483 692 523
rect 582 428 692 483
rect 582 388 617 428
rect 658 388 692 428
rect 582 368 692 388
rect 1538 501 1643 1782
rect 1538 461 1563 501
rect 1604 461 1643 501
rect 1538 412 1643 461
rect 1538 372 1563 412
rect 1604 372 1643 412
rect 242 76 347 155
rect 242 36 278 76
rect 319 36 347 76
rect -292 -354 -187 -149
rect -292 -394 -267 -354
rect -226 -394 -187 -354
rect -292 -443 -187 -394
rect -292 -483 -267 -443
rect -226 -483 -187 -443
rect -292 -617 -187 -483
rect -87 -354 26 -149
rect -87 -394 -48 -354
rect -7 -394 26 -354
rect -87 -449 26 -394
rect -87 -489 -52 -449
rect -11 -489 26 -449
rect -87 -617 26 -489
rect 242 -494 347 36
rect 242 -534 267 -494
rect 308 -534 347 -494
rect 242 -583 347 -534
rect 242 -623 267 -583
rect 308 -623 347 -583
rect 242 -757 347 -623
rect 447 -494 560 155
rect 447 -534 486 -494
rect 527 -534 560 -494
rect 447 -589 560 -534
rect 447 -629 482 -589
rect 523 -629 560 -589
rect 447 -757 560 -629
rect 1538 -411 1643 372
rect 1538 -451 1563 -411
rect 1604 -451 1643 -411
rect 1538 -500 1643 -451
rect 1538 -540 1563 -500
rect 1604 -540 1643 -500
rect 1538 -674 1643 -540
rect 1743 1911 1856 2056
rect 1743 1871 1782 1911
rect 1823 1871 1856 1911
rect 1743 1816 1856 1871
rect 1743 1776 1778 1816
rect 1819 1776 1856 1816
rect 1743 501 1856 1776
rect 1743 461 1782 501
rect 1823 461 1856 501
rect 1743 406 1856 461
rect 1743 366 1778 406
rect 1819 366 1856 406
rect 1743 -411 1856 366
rect 1743 -451 1782 -411
rect 1823 -451 1856 -411
rect 1743 -506 1856 -451
rect 1743 -546 1778 -506
rect 1819 -546 1856 -506
rect 1743 -674 1856 -546
<< pdiff >>
rect 830 2413 936 2645
rect 831 2354 936 2413
rect 831 2314 856 2354
rect 897 2314 936 2354
rect 831 2265 936 2314
rect 831 2225 856 2265
rect 897 2225 936 2265
rect 831 2124 936 2225
rect 831 2084 856 2124
rect 897 2084 936 2124
rect 831 2035 936 2084
rect 831 1995 856 2035
rect 897 1995 936 2035
rect 831 1574 936 1995
rect 831 1534 865 1574
rect 906 1534 936 1574
rect -28 1253 77 1307
rect -28 1213 5 1253
rect 46 1213 77 1253
rect -28 954 77 1213
rect -28 914 -3 954
rect 38 914 77 954
rect -28 865 77 914
rect -28 825 -3 865
rect 38 825 77 865
rect -28 691 77 825
rect 177 1242 290 1307
rect 177 1202 215 1242
rect 256 1202 290 1242
rect 177 954 290 1202
rect 177 914 216 954
rect 257 914 290 954
rect 177 859 290 914
rect 177 819 212 859
rect 253 819 290 859
rect 177 691 290 819
rect 401 1242 506 1307
rect 401 1202 437 1242
rect 478 1202 506 1242
rect 401 954 506 1202
rect 401 914 426 954
rect 467 914 506 954
rect 401 865 506 914
rect 401 825 426 865
rect 467 825 506 865
rect 401 691 506 825
rect 606 954 719 1307
rect 606 914 645 954
rect 686 914 719 954
rect 606 859 719 914
rect 606 819 641 859
rect 682 819 719 859
rect 606 691 719 819
rect 831 1073 936 1534
rect 831 1033 856 1073
rect 897 1033 936 1073
rect 831 984 936 1033
rect 831 944 856 984
rect 897 944 936 984
rect 831 810 936 944
rect 1036 2354 1149 2645
rect 1036 2314 1075 2354
rect 1116 2314 1149 2354
rect 1036 2259 1149 2314
rect 1036 2219 1071 2259
rect 1112 2219 1149 2259
rect 1036 2124 1149 2219
rect 1036 2084 1075 2124
rect 1116 2084 1149 2124
rect 1036 2029 1149 2084
rect 1036 1989 1071 2029
rect 1112 1989 1149 2029
rect 1036 1902 1149 1989
rect 1036 1862 1075 1902
rect 1116 1862 1149 1902
rect 1036 1073 1149 1862
rect 1036 1033 1075 1073
rect 1116 1033 1149 1073
rect 1036 978 1149 1033
rect 1036 938 1071 978
rect 1112 938 1149 978
rect 1036 810 1149 938
<< ndiffc >>
rect -516 1525 -489 1556
rect -516 -56 -489 -25
rect -440 1511 -413 1542
rect -440 -70 -413 -39
rect -368 1514 -341 1545
rect -368 -67 -341 -36
rect -247 1505 -220 1536
rect 1563 1871 1604 1911
rect 1563 1782 1604 1822
rect 1 483 42 523
rect 1 394 42 434
rect 220 483 261 523
rect 216 388 257 428
rect 402 483 443 523
rect 402 394 443 434
rect 621 483 662 523
rect 617 388 658 428
rect 1563 461 1604 501
rect 1563 372 1604 412
rect -248 -78 -221 -47
rect 278 36 319 76
rect -267 -394 -226 -354
rect -267 -483 -226 -443
rect -48 -394 -7 -354
rect -52 -489 -11 -449
rect 267 -534 308 -494
rect 267 -623 308 -583
rect 486 -534 527 -494
rect 482 -629 523 -589
rect 1563 -451 1604 -411
rect 1563 -540 1604 -500
rect 1782 1871 1823 1911
rect 1778 1776 1819 1816
rect 1782 461 1823 501
rect 1778 366 1819 406
rect 1782 -451 1823 -411
rect 1778 -546 1819 -506
<< pdiffc >>
rect 856 2314 897 2354
rect 856 2225 897 2265
rect 856 2084 897 2124
rect 856 1995 897 2035
rect 865 1534 906 1574
rect 5 1213 46 1253
rect -3 914 38 954
rect -3 825 38 865
rect 215 1202 256 1242
rect 216 914 257 954
rect 212 819 253 859
rect 437 1202 478 1242
rect 426 914 467 954
rect 426 825 467 865
rect 645 914 686 954
rect 641 819 682 859
rect 856 1033 897 1073
rect 856 944 897 984
rect 1075 2314 1116 2354
rect 1071 2219 1112 2259
rect 1075 2084 1116 2124
rect 1071 1989 1112 2029
rect 1075 1862 1116 1902
rect 1075 1033 1116 1073
rect 1071 938 1112 978
<< psubdiff >>
rect -184 258 -66 287
rect -184 188 -169 258
rect -99 188 -66 258
rect -184 168 -66 188
<< nsubdiff >>
rect 556 1693 594 1698
rect 527 1684 652 1693
rect 527 1654 563 1684
rect 586 1654 652 1684
rect 527 1641 652 1654
<< psubdiffcont >>
rect -169 188 -99 258
<< nsubdiffcont >>
rect 563 1654 586 1684
<< poly >>
rect 936 2645 1036 2668
rect 75 1422 188 1439
rect 75 1339 96 1422
rect 161 1339 188 1422
rect 75 1316 188 1339
rect 506 1421 606 1436
rect 506 1338 529 1421
rect 594 1338 606 1421
rect 77 1307 177 1316
rect 506 1307 606 1338
rect 1643 2056 1743 2079
rect 936 751 1036 810
rect 936 714 954 751
rect 986 714 1036 751
rect 936 697 1036 714
rect 77 645 177 691
rect 506 645 606 691
rect 81 547 181 581
rect 482 547 582 581
rect 81 309 181 368
rect 482 360 582 368
rect 81 271 99 309
rect 146 271 181 309
rect 81 247 181 271
rect 481 315 582 360
rect 481 277 512 315
rect 559 277 582 315
rect 481 248 582 277
rect 81 246 180 247
rect 347 155 447 180
rect -187 -149 -87 -101
rect -187 -632 -87 -617
rect -188 -815 -85 -632
rect 1643 -687 1743 -674
rect -188 -850 -161 -815
rect -107 -850 -85 -815
rect -188 -895 -85 -850
rect 347 -808 447 -757
rect 347 -843 367 -808
rect 421 -843 447 -808
rect 1641 -793 1743 -687
rect 1641 -826 1671 -793
rect 1719 -826 1743 -793
rect 1641 -829 1743 -826
rect 1647 -841 1741 -829
rect 347 -864 447 -843
<< polycont >>
rect 96 1339 161 1422
rect 529 1338 594 1421
rect 954 714 986 751
rect 99 271 146 309
rect 512 277 559 315
rect -161 -850 -107 -815
rect 367 -843 421 -808
rect 1671 -826 1719 -793
<< ndiffres >>
rect -521 1556 -484 1573
rect -521 1525 -516 1556
rect -489 1525 -484 1556
rect -521 -25 -484 1525
rect -521 -56 -516 -25
rect -489 -31 -484 -25
rect -445 1542 -408 1559
rect -445 1511 -440 1542
rect -413 1511 -408 1542
rect -489 -56 -485 -31
rect -521 -62 -485 -56
rect -445 -39 -408 1511
rect -445 -70 -440 -39
rect -413 -45 -408 -39
rect -373 1545 -336 1562
rect -373 1514 -368 1545
rect -341 1514 -336 1545
rect -373 -36 -336 1514
rect -413 -70 -409 -45
rect -445 -76 -409 -70
rect -373 -67 -368 -36
rect -341 -42 -336 -36
rect -252 1536 -215 1553
rect -252 1505 -247 1536
rect -220 1505 -215 1536
rect -341 -67 -337 -42
rect -373 -73 -337 -67
rect -252 -47 -215 1505
rect -252 -78 -248 -47
rect -221 -51 -215 -47
rect -221 -78 -216 -51
rect -252 -84 -216 -78
<< locali >>
rect 841 2354 907 2367
rect 841 2314 856 2354
rect 897 2314 907 2354
rect 841 2296 907 2314
rect 1061 2354 1127 2367
rect 1061 2314 1075 2354
rect 1116 2314 1127 2354
rect 1061 2296 1127 2314
rect 841 2265 907 2278
rect 841 2225 856 2265
rect 897 2225 907 2265
rect 841 2207 907 2225
rect 1061 2259 1127 2279
rect 1061 2219 1071 2259
rect 1112 2219 1127 2259
rect 1061 2208 1127 2219
rect 841 2124 907 2137
rect 841 2084 856 2124
rect 897 2084 907 2124
rect 841 2066 907 2084
rect 1061 2124 1127 2137
rect 1061 2084 1075 2124
rect 1116 2084 1127 2124
rect 1061 2066 1127 2084
rect 841 2035 907 2048
rect 841 1995 856 2035
rect 897 1995 907 2035
rect 841 1977 907 1995
rect 1061 2029 1127 2049
rect 1061 1989 1071 2029
rect 1112 1989 1127 2029
rect 1061 1978 1127 1989
rect 1065 1909 1131 1922
rect 1548 1911 1614 1924
rect 1548 1909 1563 1911
rect 1065 1902 1563 1909
rect 1065 1862 1075 1902
rect 1116 1871 1563 1902
rect 1604 1871 1614 1911
rect 1116 1869 1614 1871
rect 1116 1862 1131 1869
rect 1065 1851 1131 1862
rect 1548 1853 1614 1869
rect 1768 1911 1834 1924
rect 1768 1871 1782 1911
rect 1823 1871 1834 1911
rect 1768 1853 1834 1871
rect 1548 1822 1614 1835
rect 1548 1782 1563 1822
rect 1604 1782 1614 1822
rect 1548 1764 1614 1782
rect 1768 1816 1834 1836
rect 1768 1776 1778 1816
rect 1819 1776 1834 1816
rect 1768 1765 1834 1776
rect 549 1686 681 1693
rect 549 1684 687 1686
rect 549 1680 563 1684
rect 547 1654 563 1680
rect 586 1654 687 1684
rect 547 1628 687 1654
rect -150 1617 -112 1618
rect -522 1588 -110 1617
rect -520 1561 -482 1588
rect -150 1586 -112 1588
rect -149 1564 -112 1586
rect 651 1575 687 1628
rect 850 1575 916 1587
rect 651 1574 916 1575
rect 651 1571 865 1574
rect 35 1564 865 1571
rect -371 1562 -337 1564
rect -519 1556 -484 1561
rect -519 1525 -516 1556
rect -489 1525 -484 1556
rect -519 1522 -484 1525
rect -518 1514 -484 1522
rect -443 1559 -409 1560
rect -443 1551 -408 1559
rect -371 1551 -336 1562
rect -149 1556 865 1564
rect -236 1553 -213 1555
rect -443 1545 -336 1551
rect -443 1542 -368 1545
rect -443 1511 -440 1542
rect -413 1516 -368 1542
rect -413 1511 -408 1516
rect -371 1514 -368 1516
rect -341 1514 -336 1545
rect -249 1536 -213 1553
rect -371 1511 -336 1514
rect -443 1508 -408 1511
rect -442 1500 -408 1508
rect -370 1503 -336 1511
rect -307 1533 -279 1536
rect -250 1533 -247 1536
rect -307 1505 -247 1533
rect -220 1518 -213 1536
rect -149 1552 441 1556
rect -149 1532 217 1552
rect 244 1536 441 1552
rect 468 1536 865 1556
rect 244 1534 865 1536
rect 906 1534 916 1574
rect 244 1532 916 1534
rect -149 1521 916 1532
rect -220 1505 -215 1518
rect 850 1516 916 1521
rect -307 1501 -215 1505
rect -307 1117 -279 1501
rect -249 1494 -215 1501
rect 72 1438 193 1446
rect 72 1422 607 1438
rect 4 1382 41 1385
rect 72 1382 96 1422
rect 4 1349 96 1382
rect 4 1266 41 1349
rect 72 1339 96 1349
rect 161 1421 607 1422
rect 161 1339 529 1421
rect 72 1338 529 1339
rect 594 1338 607 1421
rect 72 1321 607 1338
rect 72 1315 193 1321
rect -9 1253 57 1266
rect -9 1213 5 1253
rect 46 1213 57 1253
rect -9 1195 57 1213
rect 201 1242 267 1255
rect 201 1202 215 1242
rect 256 1202 267 1242
rect 201 1184 267 1202
rect 423 1242 489 1255
rect 423 1202 437 1242
rect 478 1202 489 1242
rect 423 1184 489 1202
rect -307 890 -277 1117
rect 841 1073 907 1086
rect 841 1033 856 1073
rect 897 1033 907 1073
rect 841 1015 907 1033
rect 1061 1073 1127 1086
rect 1061 1033 1075 1073
rect 1116 1033 1127 1073
rect 1061 1015 1127 1033
rect 841 984 907 997
rect -18 954 48 967
rect -18 914 -3 954
rect 38 914 48 954
rect -18 896 48 914
rect 202 954 268 967
rect 202 914 216 954
rect 257 914 268 954
rect 202 896 268 914
rect 411 954 477 967
rect 411 914 426 954
rect 467 914 477 954
rect 411 896 477 914
rect 631 954 697 967
rect 631 914 645 954
rect 686 914 697 954
rect 841 944 856 984
rect 897 944 907 984
rect 841 926 907 944
rect 1061 978 1127 998
rect 1061 938 1071 978
rect 1112 938 1127 978
rect 1061 927 1127 938
rect 631 896 697 914
rect -305 859 -277 890
rect 1071 887 1104 927
rect -309 804 -277 859
rect -18 865 48 878
rect -18 825 -3 865
rect 38 825 48 865
rect -18 807 48 825
rect 202 859 268 879
rect 202 819 212 859
rect 253 819 268 859
rect 202 808 268 819
rect 411 865 477 878
rect 411 825 426 865
rect 467 825 477 865
rect 631 859 697 879
rect 631 846 641 859
rect 411 807 477 825
rect 628 819 641 846
rect 682 819 697 859
rect 628 808 697 819
rect 1071 846 1365 887
rect 1071 813 1104 846
rect -309 368 -278 804
rect 5 536 32 807
rect 628 602 673 808
rect 1056 757 1098 771
rect 944 751 1098 757
rect 944 714 954 751
rect 986 714 1098 751
rect 944 710 1098 714
rect 1056 622 1098 710
rect 1056 602 1080 622
rect 1170 602 1200 846
rect 628 563 1080 602
rect 1152 594 1231 602
rect 1152 567 1205 594
rect 1228 567 1231 594
rect 1152 563 1231 567
rect 628 536 673 563
rect -14 523 52 536
rect -14 483 1 523
rect 42 483 52 523
rect -14 465 52 483
rect 206 523 272 536
rect 206 483 220 523
rect 261 483 272 523
rect 206 465 272 483
rect 387 523 453 536
rect 387 483 402 523
rect 443 483 453 523
rect 387 465 453 483
rect 607 523 673 536
rect 607 483 621 523
rect 662 483 673 523
rect 607 465 673 483
rect 1548 501 1614 514
rect 1548 461 1563 501
rect 1604 461 1614 501
rect -14 434 52 447
rect -14 394 1 434
rect 42 394 52 434
rect -14 376 52 394
rect 206 430 272 448
rect 387 434 453 447
rect 387 430 402 434
rect 206 428 402 430
rect 206 388 216 428
rect 257 394 402 428
rect 443 394 453 434
rect 257 388 453 394
rect 206 382 453 388
rect 206 377 272 382
rect -530 -25 -476 -11
rect -530 -56 -516 -25
rect -489 -47 -476 -25
rect -454 -39 -400 -25
rect -454 -47 -440 -39
rect -489 -56 -440 -47
rect -530 -69 -440 -56
rect -530 -85 -481 -69
rect -454 -70 -440 -69
rect -413 -70 -400 -39
rect -454 -74 -400 -70
rect -382 -36 -328 -22
rect -382 -67 -368 -36
rect -341 -67 -328 -36
rect -382 -71 -328 -67
rect -451 -82 -400 -74
rect -379 -83 -328 -71
rect -310 -83 -278 368
rect 213 332 256 377
rect 387 376 453 382
rect 607 428 673 448
rect 1548 443 1614 461
rect 1768 501 1834 514
rect 1768 461 1782 501
rect 1823 461 1834 501
rect 1768 443 1834 461
rect 607 388 617 428
rect 658 388 673 428
rect 607 377 673 388
rect 1548 412 1614 425
rect 1548 372 1563 412
rect 1604 372 1614 412
rect 1548 354 1614 372
rect 1768 406 1834 426
rect 1768 366 1778 406
rect 1819 366 1834 406
rect 1768 355 1834 366
rect 87 309 166 325
rect 87 271 99 309
rect 146 271 166 309
rect -182 258 -34 266
rect -182 188 -169 258
rect -99 188 -34 258
rect -182 177 -34 188
rect 87 225 166 271
rect 87 187 102 225
rect 149 187 166 225
rect 87 182 166 187
rect 210 214 256 332
rect 494 315 573 333
rect 494 277 512 315
rect 559 277 573 315
rect 494 236 573 277
rect 274 214 328 216
rect 210 186 328 214
rect 494 198 508 236
rect 555 198 573 236
rect 494 190 573 198
rect 216 180 328 186
rect 274 89 328 180
rect 263 76 329 89
rect 263 36 278 76
rect 319 36 329 76
rect -254 -47 -215 -39
rect -254 -78 -248 -47
rect -221 -73 -215 -47
rect -221 -74 -214 -73
rect -221 -78 -212 -74
rect -254 -83 -212 -78
rect -379 -95 -278 -83
rect -379 -108 -279 -95
rect -256 -106 -212 -83
rect -373 -111 -279 -108
rect -369 -112 -346 -111
rect -249 -142 -214 -106
rect -248 -198 -216 -142
rect -270 -269 -204 -198
rect 263 -313 329 36
rect -282 -354 -216 -341
rect -282 -394 -267 -354
rect -226 -394 -216 -354
rect -282 -412 -216 -394
rect -62 -354 4 -341
rect -62 -394 -48 -354
rect -7 -394 4 -354
rect -62 -412 4 -394
rect 1548 -411 1614 -398
rect -282 -443 -216 -430
rect -282 -483 -267 -443
rect -226 -483 -216 -443
rect -282 -501 -216 -483
rect -62 -449 4 -429
rect -62 -489 -52 -449
rect -11 -489 4 -449
rect 1548 -451 1563 -411
rect 1604 -451 1614 -411
rect 1548 -469 1614 -451
rect 1768 -411 1834 -398
rect 1768 -451 1782 -411
rect 1823 -451 1834 -411
rect 1768 -469 1834 -451
rect -62 -500 4 -489
rect 252 -494 318 -481
rect -272 -815 -230 -501
rect 252 -534 267 -494
rect 308 -534 318 -494
rect 252 -552 318 -534
rect 472 -494 538 -481
rect 472 -534 486 -494
rect 527 -534 538 -494
rect 472 -552 538 -534
rect 1548 -500 1614 -487
rect 1548 -540 1563 -500
rect 1604 -540 1614 -500
rect 1548 -558 1614 -540
rect 1768 -506 1834 -486
rect 1768 -546 1778 -506
rect 1819 -546 1834 -506
rect 1768 -557 1834 -546
rect 252 -583 318 -570
rect 252 -623 267 -583
rect 308 -623 318 -583
rect 252 -641 318 -623
rect 472 -589 538 -569
rect 472 -629 482 -589
rect 523 -629 538 -589
rect 472 -636 489 -629
rect 507 -636 538 -629
rect 472 -640 538 -636
rect 342 -792 1755 -775
rect -176 -793 1755 -792
rect -176 -808 1671 -793
rect -176 -815 367 -808
rect -290 -850 -161 -815
rect -107 -843 367 -815
rect 421 -826 1671 -808
rect 1719 -826 1755 -793
rect 421 -843 1755 -826
rect -107 -846 1755 -843
rect -107 -850 436 -846
rect -290 -862 436 -850
rect -176 -868 436 -862
rect 1788 -942 1811 -557
rect 1701 -981 1811 -942
rect -135 -984 1811 -981
rect -135 -1023 -45 -984
rect -23 -996 1811 -984
rect -23 -1023 492 -996
rect 509 -1023 1811 -996
rect -135 -1040 1811 -1023
<< viali >>
rect 217 1532 244 1552
rect 441 1536 468 1556
rect 219 1216 247 1238
rect 441 1216 469 1238
rect 1205 567 1228 594
rect 102 187 149 225
rect 508 198 555 236
rect -42 -488 -23 -466
rect 489 -629 507 -607
rect 489 -636 507 -629
rect -45 -1023 -23 -984
rect 492 -1023 509 -996
<< metal1 >>
rect 212 1552 254 1561
rect 212 1532 217 1552
rect 244 1532 254 1552
rect 212 1238 254 1532
rect 212 1216 219 1238
rect 247 1216 254 1238
rect 212 1209 254 1216
rect 434 1556 476 1561
rect 434 1536 441 1556
rect 468 1536 476 1556
rect 434 1238 476 1536
rect 434 1216 441 1238
rect 469 1216 476 1238
rect 434 1209 476 1216
rect 1198 594 1264 602
rect 1198 567 1205 594
rect 1228 567 1264 594
rect 1198 563 1264 567
rect 504 236 561 242
rect 98 225 155 233
rect 98 187 102 225
rect 149 187 155 225
rect 98 168 155 187
rect 504 198 508 236
rect 555 205 561 236
rect 555 198 741 205
rect 504 177 741 198
rect 507 172 741 177
rect -50 -466 -15 -455
rect -50 -488 -42 -466
rect -23 -488 -15 -466
rect -50 -984 -15 -488
rect -50 -1023 -45 -984
rect -23 -1023 -15 -984
rect -50 -1040 -15 -1023
rect 485 -607 514 -599
rect 485 -636 489 -607
rect 507 -636 514 -607
rect 485 -996 514 -636
rect 485 -1023 492 -996
rect 509 -1023 514 -996
rect 485 -1031 514 -1023
<< labels >>
rlabel locali 64 1534 64 1534 1 vdd
rlabel metal1 1247 579 1247 579 1 out2
rlabel metal1 121 174 121 174 1 in1
rlabel metal1 688 188 688 188 1 in2
rlabel locali -54 212 -54 212 1 vss
rlabel locali 815 -1015 815 -1015 1 vss
<< end >>
