magic
tech sky130A
timestamp 1651363021
<< metal3 >>
rect 1485 6163 5441 6164
rect 556 5985 5441 6163
rect 556 5896 5436 5985
rect 1409 5893 5436 5896
rect 536 3161 643 3177
rect -6674 3123 -5651 3126
rect -1482 3123 643 3161
rect -6674 2947 643 3123
rect -6674 2933 -5498 2947
rect -1482 2946 643 2947
rect -6674 2839 -5651 2933
rect 536 2897 643 2946
rect -9482 1657 -7891 1660
rect -9482 1652 -6574 1657
rect -10398 1644 -6574 1652
rect -11675 1514 -6574 1644
rect -11675 1346 -9378 1514
rect -8091 1512 -6574 1514
rect -10398 1343 -9378 1346
<< metal4 >>
rect -11219 -115 -11110 286
rect -9934 -61 -9845 275
rect -8616 -67 -8521 235
rect -6214 -51 -6119 251
rect -3606 50 -3489 395
rect 4242 -73 4359 272
use mimcap1C  mimcap1C_1
timestamp 1649877290
transform 1 0 -11460 0 1 567
box -220 -375 810 905
use mimcap1C  mimcap1C_0
timestamp 1649877290
transform 1 0 -10185 0 1 542
box -220 -375 810 905
use mimcap2C  mimcap2C_0
timestamp 1649877975
transform 1 0 -9074 0 1 279
box 0 -100 2115 1380
use mimcap4C  mimcap4C_0
timestamp 1650135350
transform 1 0 -6683 0 1 1561
box 0 -1395 2120 1480
use mimcap8C  mimcap8C_0
timestamp 1651320701
transform 1 0 -4067 0 1 219
box 0 -100 4290 2975
use mimcap16C  mimcap16C_0
timestamp 1651320701
transform -1 0 4835 0 1 3123
box 0 -2990 4300 3075
<< labels >>
rlabel metal3 5124 6041 5124 6041 1 vcommon
rlabel metal4 -8594 -33 -8594 -33 1 C2
rlabel metal4 -6184 -30 -6184 -30 1 C4
rlabel metal4 -3560 84 -3560 84 1 C8
rlabel metal4 4242 -73 4359 272 1 C16
rlabel metal4 -9896 -16 -9896 -16 1 C1
rlabel metal4 -11188 -18 -11188 -18 1 C0
<< end >>
