** sch_path: /home/rperry/saradcspr2022/top.sch


.param vONE=2
.param vadc=1.5


**.subckt top dataOut[2] dataOut[1] dataOut[0] nEndCnv
*.opin dataOut[2]
*.opin dataOut[1]
*.opin dataOut[0]
*.opin nEndCnv
x1 CompOut SH VREF B0 B1 B2 AGND dacVin dacblock
x2 dacVin Vin SH ug_sample_hold
Vmax VDD GND 2
Vmax1 Vin GND sin(1.5 0.5 10000 2u )
Vmax3 AGND GND 1
Vmax4 VREF GND 2
x3 GND VDD reset clock nStartCnv SH B2 B1 B0 CompOut dataOut[2] dataOut[1] dataOut[0] nEndCnv
+ sar3bitsreg
V4 reset GND DC 0 pwl (0n 0 500n 0 510n 2)
V1 clock GND DC 2 pulse(0 2 0 10n 10n 1u 2u)
V3 nStartCnv GND dc 2 pwl (0n 2 1.5u 2 1.51u 0)
**** begin user architecture code


.include ./spice/opamp_sky130.sp
.include ./spice/sar3bitsreg.sp

.op
.control
run
**plot i(Vswitch)

.endc



** opencircuitdesign pdks install
.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.include /usr/local/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice
.include /usr/local/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_ef_sc_hd__decap_12.spice



**** end user architecture code
**.ends

* expanding   symbol:  dacblock.sym # of pins=8
** sym_path: /home/rperry/saradcspr2022/dacblock.sym
** sch_path: /home/rperry/saradcspr2022/dacblock.sch
.subckt dacblock  CompOut SH VREF B0 B1 B2 AGND Vin
*.ipin Vin
*.ipin AGND
*.ipin VREF
*.ipin SH
*.ipin B0
*.ipin B1
*.ipin B2
*.opin CompOut
XC1 Vcommon c1v sky130_fd_pr__cap_mim_m3_1 W=10 L=10 MF=1 m=1
XC2 Vcommon c2v sky130_fd_pr__cap_mim_m3_1 W=10 L=10 MF=1 m=1
x3 Vcommon AGND CompOut skywater_comparator
XC6 Vcommon c4v sky130_fd_pr__cap_mim_m3_1 W=10 L=10 MF=4 m=4
XC7 Vcommon c3v sky130_fd_pr__cap_mim_m3_1 W=10 L=10 MF=2 m=2
x1 c4v SH Vin AGND VREF AGND B2 4x1analogmux
x2 c3v SH Vin AGND VREF AGND B1 4x1analogmux
x4 c2v SH Vin AGND VREF AGND B0 4x1analogmux
x5 c1v Vin AGND SH 2x1analogmux
x6 AGND SH Vcommon analog_switch
.ends


* expanding   symbol:  ug_sample_hold.sym # of pins=3
** sym_path: /home/rperry/saradcspr2022/ug_sample_hold.sym
** sch_path: /home/rperry/saradcspr2022/ug_sample_hold.sch
.subckt ug_sample_hold  Vout Vin SHClk
*.ipin Vin
*.ipin SHClk
*.opin Vout
x1 Vin SHClk Vout analog_switch
.ends


* expanding   symbol:  skywater_comparator.sym # of pins=3
** sym_path: /home/rperry/saradcspr2022/skywater_comparator.sym
** sch_path: /home/rperry/saradcspr2022/skywater_comparator.sch
.subckt skywater_comparator  Vmin Vpos Y
*.ipin Vpos
*.ipin Vmin
*.opin Y
x1 Y net1 VDD GND not W_N=1 L_N=0.15 W_P=2 L_P=0.15 m=10
x2 Vmin Vpos net1 VDD GND opamp_sky130
.ends


* expanding   symbol:  4x1analogmux.sym # of pins=7
** sym_path: /home/rperry/saradcspr2022/4x1analogmux.sym
** sch_path: /home/rperry/saradcspr2022/4x1analogmux.sch
.subckt 4x1analogmux  Vout S1 A3 A2 A1 A0 S0
*.ipin A3
*.ipin A2
*.ipin A1
*.ipin A0
*.ipin S1
*.ipin S0
*.opin Vout
x2 net2 A1 A0 S0 2x1analogmux
x3 Vout net1 net2 S1 2x1analogmux
x1 net1 A3 A2 S0 2x1analogmux
.ends


* expanding   symbol:  2x1analogmux.sym # of pins=4
** sym_path: /home/rperry/saradcspr2022/2x1analogmux.sym
** sch_path: /home/rperry/saradcspr2022/2x1analogmux.sch
.subckt 2x1analogmux  Vout A1 A0 S
*.ipin S
*.opin Vout
*.ipin A1
*.ipin A0
x1 net1 A1 Vout S dacpassgate
x2 S A0 Vout net1 dacpassgate
x3 net1 S VDD GND not W_N=1 L_N=0.15 W_P=2 L_P=0.15 m=1
.ends


* expanding   symbol:  analog_switch.sym # of pins=3
** sym_path: /home/rperry/saradcspr2022/analog_switch.sym
** sch_path: /home/rperry/saradcspr2022/analog_switch.sch
.subckt analog_switch  Vin S Vout
*.ipin S
*.ipin Vin
*.opin Vout
x1 net1 Vin Vout S dacpassgate
x2 net1 S VDD GND not W_N=1 L_N=0.15 W_P=2 L_P=0.15 m=1
.ends


* expanding   symbol:  not.sym # of pins=2
** sym_path: /home/rperry/saradcspr2022/not.sym
** sch_path: /home/rperry/saradcspr2022/not.sch
.subckt not  y a  VCCPIN  VSSPIN      W_N=1 L_N=0.15 W_P=2 L_P=0.15
*.opin y
*.ipin a
XM1 y a VSSPIN VSSPIN sky130_fd_pr__nfet_01v8 L=L_N W=W_N nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 y a VCCPIN VCCPIN sky130_fd_pr__pfet_01v8 L=L_P W=W_P nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  dacpassgate.sym # of pins=4
** sym_path: /home/rperry/saradcspr2022/dacpassgate.sym
** sch_path: /home/rperry/saradcspr2022/dacpassgate.sch
.subckt dacpassgate  GP A Z GN
*.iopin A
*.iopin Z
*.ipin GP
*.ipin GN
XM1 Z GN A GND sky130_fd_pr__nfet_01v8 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=10 m=10
XM2 Z GP A VDD sky130_fd_pr__pfet_01v8 L=0.5 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=10 m=10
.ends

.GLOBAL GND
.GLOBAL VDD
.end
