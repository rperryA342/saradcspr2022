** sch_path: /home/reg/saradcspr2022/dac5bitsblock_test.sch


.param vONE=2
.param AGND=1
.param rt=5n
.param pw=10u
.param t0=100n
.param t0r=t0+rt
.param t1=t0r+pw
.param t1r=t1+rt
.param t2=t1r+pw
.param t2r=t2+rt
.param t3=t2r+pw
.param t3r=t3+rt
.param t4=t3r+pw
.param t4r=t4+rt
.param t5=t4r+pw
.param t5r=t5+rt
.param t6=t5r+pw
.param t6r=t6+rt
.param t7=t6r+pw
.param t7r=t7+rt
.param t8=t7r+pw
.param t8r=t8+rt
.param t9=t8r+pw
.param t9r=t9+rt
.param t10=t9r+pw
.param t10r=t10+rt
.param t11=t10r+pw
.param t11r=t11+rt

.param b4d=VONE
.param b3d=0
.param b2d=VONE
.param b1d=0
.param b0d=VONE
.param vpcomp=(b4d/2)+(b3d/4)+(b2d/8)+(b1d/16)+(b0d/32)
.param vadc=(vpcomp/2)+AGND



**.subckt dac5bitsblock_test
Vmax VDD GND 2
Vmax1 Vin GND {vadc}
Vmax3 AGND GND 1
V4 SH GND DC 0 pwl (0n 0 {t0} 0 {t0r} 2 {t1} 2 {t1r} 0)
Vmax4 VREF GND 2
V1 B3 GND DC 0 pwl (0n 0 {t0} 0 {t0r} 2 {t1} 2 {t1r} 0 {t4} 0 {t4r} 2 {t5} 2 {t5r} {b3d})
V3 B2 GND dc 0 pwl (0n 0 {t0} 0 {t0r} 2 {t1} 2 {t1r} 0 {t6} 0 {t6r} 2 {t7} 2 {t7r} {b2d})
V5 B4 GND DC 0 pwl (0n 0 {t0} 0 {t0r} 2 {t1} 2 {t1r} 0 {t2} 0 {t2r} 2 {t3} 2 {t3r} {b4d})
XC3 AGND GND sky130_fd_pr__cap_mim_m3_1 W=10 L=10 MF=1 m=1
x1 CompOut SH VREF B4 B3 B2 B1 B0 AGND Vin dacblock5bits
V2 B1 GND DC 0 pwl (0n 0 {t0} 0 {t0r} 2 {t1} 2 {t1r} 0 {t8} 0 {t8r} 2 {t9} 2 {t9r} {b1d})
V6 B0 GND DC 0 pwl (0n 0 {t0} 0 {t0r} 2 {t1} 2 {t1r} 0 {t10} 0 {t10r} 2 {t11} 2 {t11r} {b0d})
C1 CompOut GND 1p m=1
**** begin user architecture code


**.include spice/caparray.sp

.tran 0.1u 120u
.control
run
plot v(CompOut) v(x1.vcommon)

.endc



** opencircuitdesign pdks install
.lib /home/reg/OpenLane/pdks/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.include /home/reg/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice
.include /home/reg/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_ef_sc_hd__decap_12.spice



**** end user architecture code
**.ends

* expanding   symbol:  dacblock5bits.sym # of pins=10
** sym_path: /home/reg/saradcspr2022/dacblock5bits.sym
** sch_path: /home/reg/saradcspr2022/dacblock5bits.sch
.subckt dacblock5bits  CompOut SH VREF B4 B3 B2 B1 B0 AGND Vin
*.ipin B0
*.ipin B1
*.ipin B2
*.ipin B3
*.ipin B4
*.ipin Vin
*.ipin SH
*.opin CompOut
*.iopin AGND
*.iopin VREF
x1 C16 SH Vin AGND VREF AGND B4 4x1analogmux
x2 C8 SH Vin AGND VREF AGND B3 4x1analogmux
x4 C4 SH Vin AGND VREF AGND B2 4x1analogmux
x5 C0 Vin AGND SH 2x1analogmux
x6 AGND SH vcommon analog_switch
x7 C2 SH Vin AGND VREF AGND B1 4x1analogmux
x8 C1 SH Vin AGND VREF AGND B0 4x1analogmux
x9 vcommon C0 C1 C2 C4 C8 C16 caparray
x3 AGND vcommon CompOut VDD GND simpleComp
.ends


* expanding   symbol:  4x1analogmux.sym # of pins=7
** sym_path: /home/reg/saradcspr2022/4x1analogmux.sym
** sch_path: /home/reg/saradcspr2022/4x1analogmux.sch
.subckt 4x1analogmux  Vout S1 A3 A2 A1 A0 S0
*.ipin A3
*.ipin A2
*.ipin A1
*.ipin A0
*.ipin S1
*.ipin S0
*.opin Vout
x2 nS1S0 A1 A0 S0 2x1analogmux
x3 Vout S1S0 nS1S0 S1 2x1analogmux
x1 S1S0 A3 A2 S0 2x1analogmux
.ends


* expanding   symbol:  2x1analogmux.sym # of pins=4
** sym_path: /home/reg/saradcspr2022/2x1analogmux.sym
** sch_path: /home/reg/saradcspr2022/2x1analogmux.sch
.subckt 2x1analogmux  Vout A1 A0 S
*.ipin S
*.opin Vout
*.ipin A1
*.ipin A0
x1 nS A1 Vout S dacpassgate
x2 S A0 Vout nS dacpassgate
x3 nS S VDD GND not W_N=1 L_N=0.15 W_P=2 L_P=0.15 m=1
.ends


* expanding   symbol:  analog_switch.sym # of pins=3
** sym_path: /home/reg/saradcspr2022/analog_switch.sym
** sch_path: /home/reg/saradcspr2022/analog_switch.sch
.subckt analog_switch  Vin S Vout
*.ipin S
*.ipin Vin
*.opin Vout
x1 nS Vin Vout S dacpassgate
x2 nS S VDD GND not W_N=1 L_N=0.15 W_P=2 L_P=0.15 m=1
.ends


* expanding   symbol:  caparray.sym # of pins=7
** sym_path: /home/reg/saradcspr2022/caparray.sym
** sch_path: /home/reg/saradcspr2022/caparray.sch
.subckt caparray  vcommon  C0  C1  C2  C4  C8  C16
*.iopin C0
*.iopin C1
*.iopin C2
*.iopin C4
*.iopin C8
*.iopin C16
*.iopin vcommon
XC1 C0 vcommon sky130_fd_pr__cap_mim_m3_1 W=100 L=100 MF=1 m=1
XC2 C1 vcommon sky130_fd_pr__cap_mim_m3_1 W=100 L=100 MF=1 m=1
XC3 C2 vcommon sky130_fd_pr__cap_mim_m3_1 W=100 L=100 MF=2 m=2
XC4 C4 vcommon sky130_fd_pr__cap_mim_m3_1 W=100 L=100 MF=4 m=4
XC5 C8 vcommon sky130_fd_pr__cap_mim_m3_1 W=100 L=100 MF=8 m=8
XC6 C16 vcommon sky130_fd_pr__cap_mim_m3_1 W=100 L=100 MF=16 m=16
.ends


* expanding   symbol:  simpleComp.sym # of pins=5
** sym_path: /home/reg/saradcspr2022/simpleComp.sym
** sch_path: /home/reg/saradcspr2022/simpleComp.sch
.subckt simpleComp  Vm Vp Vout VDDPIN GNDPIN
*.ipin Vp
*.ipin Vm
*.opin Vout
*.iopin VDDPIN
*.iopin GNDPIN
C7 GP 0 4f m=1
XM4 SP GNDPIN VDDPIN VDDPIN sky130_fd_pr__pfet_01v8 L=1 W=0.55 nf=1 ad='W * 0.29' as='W * 0.29' pd='W + 2 * 0.29'
+ ps='W + 2 * 0.29' nrd=0 nrs=0 sa=0 sb=0 sd=0 mult=1 m=1
XM18 diffout GP GNDPIN GNDPIN sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='W * 0.29' as='W * 0.29' pd='2*(W + 0.29)'
+ ps='2*(W + 0.29)' nrd=0 nrs=0 sa=0 sb=0 sd=0 mult=1 m=1
XM19 GP GP GNDPIN GNDPIN sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='W * 0.29' as='W * 0.29' pd='2*(W + 0.29)'
+ ps='2*(W + 0.29)' nrd=0 nrs=0 sa=0 sb=0 sd=0 mult=1 m=1
XM20 diffout Vp SP VDDPIN sky130_fd_pr__pfet_01v8_lvt L=0.35 W=1 nf=1 ad='W * 0.29' as='W * 0.29' pd='2*(W + 0.29)'
+ ps='2*(W + 0.29)' nrd=0 nrs=0 sa=0 sb=0 sd=0 mult=1 m=1
XM21 GP Vm SP VDDPIN sky130_fd_pr__pfet_01v8_lvt L=0.35 W=1 nf=1 ad='W * 0.29' as='W * 0.29' pd='2*(W + 0.29)'
+ ps='2*(W + 0.29)' nrd=0 nrs=0 sa=0 sb=0 sd=0 mult=1 m=1
x1 Vout diffout VDDPIN GNDPIN not W_N=1 L_N=0.15 W_P=2 L_P=0.15 m=10
.ends


* expanding   symbol:  dacpassgate.sym # of pins=4
** sym_path: /home/reg/saradcspr2022/dacpassgate.sym
** sch_path: /home/reg/saradcspr2022/dacpassgate.sch
.subckt dacpassgate  GP A Z GN
*.iopin A
*.iopin Z
*.ipin GP
*.ipin GN
XM1 Z GN A GND sky130_fd_pr__nfet_01v8 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=10 m=10
XM2 Z GP A VDD sky130_fd_pr__pfet_01v8 L=0.5 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=10 m=10
.ends


* expanding   symbol:  not.sym # of pins=2
** sym_path: /home/reg/saradcspr2022/not.sym
** sch_path: /home/reg/saradcspr2022/not.sch
.subckt not  y a  VCCPIN  VSSPIN      W_N=1 L_N=0.15 W_P=2 L_P=0.15
*.opin y
*.ipin a
XM1 y a VSSPIN VSSPIN sky130_fd_pr__nfet_01v8 L=L_N W=W_N nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 y a VCCPIN VCCPIN sky130_fd_pr__pfet_01v8 L=L_P W=W_P nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL GND
.GLOBAL VDD
.end
