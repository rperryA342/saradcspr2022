* SPICE3 file created from caparry.ext - technology: sky130A

*.option scale=10000u

.subckt caparray vcommon B5 B0 B1 B2 B3 B4 

X50 B5 vcommon sky130_fd_pr__cap_mim_m3_1 l=100 w=100
X0  B0 vcommon sky130_fd_pr__cap_mim_m3_1 l=100 w=100
X1  B2 vcommon sky130_fd_pr__cap_mim_m3_1 l=100 w=100
X2  B2 vcommon sky130_fd_pr__cap_mim_m3_1 l=100 w=100
X3  B2 vcommon sky130_fd_pr__cap_mim_m3_1 l=100 w=100
X4  B2 vcommon sky130_fd_pr__cap_mim_m3_1 l=100 w=100
X5  B1 vcommon sky130_fd_pr__cap_mim_m3_1 l=100 w=100
X6  B1 vcommon sky130_fd_pr__cap_mim_m3_1 l=100 w=100
X7  B3 vcommon sky130_fd_pr__cap_mim_m3_1 l=100 w=100
X8  B3 vcommon sky130_fd_pr__cap_mim_m3_1 l=100 w=100
X9  B3 vcommon sky130_fd_pr__cap_mim_m3_1 l=100 w=100
X10 B3 vcommon sky130_fd_pr__cap_mim_m3_1 l=100 w=100
X11 B3 vcommon sky130_fd_pr__cap_mim_m3_1 l=100 w=100
X12 B3 vcommon sky130_fd_pr__cap_mim_m3_1 l=100 w=100
X13 B3 vcommon sky130_fd_pr__cap_mim_m3_1 l=100 w=100
X14 B3 vcommon sky130_fd_pr__cap_mim_m3_1 l=100 w=100
X15 B4 vcommon sky130_fd_pr__cap_mim_m3_1 l=100 w=100
X16 B4 vcommon sky130_fd_pr__cap_mim_m3_1 l=100 w=100
X17 B4 vcommon sky130_fd_pr__cap_mim_m3_1 l=100 w=100
X18 B4 vcommon sky130_fd_pr__cap_mim_m3_1 l=100 w=100
X19 B4 vcommon sky130_fd_pr__cap_mim_m3_1 l=100 w=100
X20 B4 vcommon sky130_fd_pr__cap_mim_m3_1 l=100 w=100
X21 B4 vcommon sky130_fd_pr__cap_mim_m3_1 l=100 w=100
X22 B4 vcommon sky130_fd_pr__cap_mim_m3_1 l=100 w=100
X23 B4 vcommon sky130_fd_pr__cap_mim_m3_1 l=100 w=100
X24 B4 vcommon sky130_fd_pr__cap_mim_m3_1 l=100 w=100
X25 B4 vcommon sky130_fd_pr__cap_mim_m3_1 l=100 w=100
X26 B4 vcommon sky130_fd_pr__cap_mim_m3_1 l=100 w=100
X27 B4 vcommon sky130_fd_pr__cap_mim_m3_1 l=100 w=100
X28 B4 vcommon sky130_fd_pr__cap_mim_m3_1 l=100 w=100
X29 B4 vcommon sky130_fd_pr__cap_mim_m3_1 l=100 w=100
X30 B4 vcommon sky130_fd_pr__cap_mim_m3_1 l=100 w=100

.ends
